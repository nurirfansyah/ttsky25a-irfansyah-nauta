magic
tech sky130A
magscale 1 2
timestamp 1757958777
<< nwell >>
rect 1200 -970 1680 360
<< pwell >>
rect 1210 -1700 1660 -1550
<< locali >>
rect 1200 330 1680 350
rect 1200 290 1230 330
rect 1650 290 1680 330
rect 1200 270 1680 290
rect 1280 -390 1590 -250
rect 1190 -2160 1670 -2140
rect 1190 -2220 1210 -2160
rect 1650 -2220 1670 -2160
rect 1190 -2240 1670 -2220
<< viali >>
rect 1230 290 1650 330
rect 1210 -2220 1650 -2160
<< metal1 >>
rect 1200 330 1680 520
rect 1200 290 1230 330
rect 1650 290 1680 330
rect 1200 270 1680 290
rect 1310 0 1360 270
rect 1400 160 1470 220
rect 980 -120 1180 -60
rect 980 -190 1470 -120
rect 980 -260 1180 -190
rect 1510 -290 1570 50
rect 1300 -350 1570 -290
rect 1300 -650 1360 -350
rect 1400 -500 1470 -440
rect 1000 -990 1200 -920
rect 1400 -990 1470 -770
rect 1000 -1070 1470 -990
rect 1000 -1120 1200 -1070
rect 1400 -1260 1470 -1070
rect 1510 -990 1550 -640
rect 1660 -990 1860 -920
rect 1510 -1070 1860 -990
rect 1000 -1660 1200 -1530
rect 1310 -1550 1360 -1320
rect 1510 -1390 1550 -1070
rect 1660 -1120 1860 -1070
rect 1400 -1470 1470 -1420
rect 1310 -1600 1560 -1550
rect 1000 -1730 1470 -1660
rect 1400 -1870 1470 -1730
rect 1310 -2140 1370 -1930
rect 1510 -1960 1560 -1600
rect 1400 -2080 1470 -2030
rect 1190 -2160 1670 -2140
rect 1190 -2220 1210 -2160
rect 1650 -2220 1670 -2160
rect 1190 -2390 1670 -2220
use sky130_fd_pr__nfet_01v8_SALLWN  XM1
timestamp 1757956269
transform 1 0 1436 0 1 -1340
box -226 -260 226 260
use sky130_fd_pr__pfet_01v8_6QYSWZ  XM2
timestamp 1757956269
transform 1 0 1436 0 1 -641
box -226 -319 226 319
use sky130_fd_pr__pfet_01v8_6QYSWZ  XM3
timestamp 1757956269
transform 1 0 1436 0 1 9
box -226 -319 226 319
use sky130_fd_pr__nfet_01v8_SALLWN  XM4
timestamp 1757956269
transform 1 0 1446 0 1 -1950
box -226 -260 226 260
<< labels >>
flabel metal1 1200 320 1400 520 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 1190 -2390 1390 -2190 0 FreeSans 256 0 0 0 gnd
port 5 nsew
flabel metal1 980 -260 1180 -60 0 FreeSans 256 0 0 0 sw_p
port 3 nsew
flabel metal1 1000 -1120 1200 -920 0 FreeSans 256 0 0 0 in
port 2 nsew
flabel metal1 1660 -1120 1860 -920 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 1000 -1730 1200 -1530 0 FreeSans 256 0 0 0 sw_n
port 4 nsew
<< end >>
