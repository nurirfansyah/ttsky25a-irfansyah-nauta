magic
tech sky130A
timestamp 1757957364
<< checkpaint >>
rect -630 190 1450 1145
rect -630 100 2100 190
rect -630 -430 2810 100
rect -630 -3230 4540 -430
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
rect 0 -1200 100 -1100
rect 0 -1400 100 -1300
rect 0 -1600 100 -1500
rect 0 -1800 100 -1700
rect 0 -2000 100 -1900
rect 0 -2200 100 -2100
rect 0 -2400 100 -2300
rect 0 -2600 100 -2500
use ff_inv  x1
timestamp 1757952934
transform 1 0 -1155 0 1 -1405
box 1155 -1195 1565 1920
use ff_inv  x2
timestamp 1757952934
transform 1 0 -745 0 1 -1405
box 1155 -1195 1565 1920
use sc_inv  x3
timestamp 1757954003
transform 1 0 270 0 1 -1325
box 550 -1275 875 885
use sc_inv  x4
timestamp 1757954003
transform 1 0 595 0 1 -1325
box 550 -1275 875 885
use cc_inv_4  x5
timestamp 1757954784
transform 1 0 1085 0 1 -1505
box 385 -1095 740 975
use cc_inv_4  x6
timestamp 1757954784
transform 1 0 1440 0 1 -1505
box 385 -1095 740 975
use cc_inv_dt05  x7
timestamp 1757956456
transform 1 0 1690 0 1 -1405
box 490 -1195 930 260
use cc_inv_dt05  x8
timestamp 1757956456
transform 1 0 2130 0 1 -1405
box 490 -1195 930 260
use cc_inv_dt05_long  x11
timestamp 1757957181
transform 1 0 2585 0 1 -1510
box 475 -1090 900 450
use cc_inv_dt05_long  x12
timestamp 1757957181
transform 1 0 3010 0 1 -1510
box 475 -1090 900 450
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 vdd
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 out_n
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 in_p
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 out_p
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 in_n
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 sw_p_A1
port 5 nsew
flabel metal1 0 -1200 100 -1100 0 FreeSans 128 0 0 0 sw_p_B1
port 6 nsew
flabel metal1 0 -1400 100 -1300 0 FreeSans 128 0 0 0 sw_p_A05
port 7 nsew
flabel metal1 0 -1600 100 -1500 0 FreeSans 128 0 0 0 sw_p_B05
port 8 nsew
flabel metal1 0 -1800 100 -1700 0 FreeSans 128 0 0 0 sw_n_A1
port 9 nsew
flabel metal1 0 -2000 100 -1900 0 FreeSans 128 0 0 0 sw_n_B1
port 10 nsew
flabel metal1 0 -2200 100 -2100 0 FreeSans 128 0 0 0 sw_n_A05
port 11 nsew
flabel metal1 0 -2400 100 -2300 0 FreeSans 128 0 0 0 sw_n_B05
port 12 nsew
flabel metal1 0 -2600 100 -2500 0 FreeSans 128 0 0 0 gnd
port 13 nsew
<< end >>
