magic
tech sky130A
magscale 1 2
timestamp 1757947919
<< error_p >>
rect -88 472 -30 478
rect 30 472 88 478
rect -88 438 -76 472
rect 30 438 42 472
rect -88 432 -30 438
rect 30 432 88 438
rect -88 -438 -30 -432
rect 30 -438 88 -432
rect -88 -472 -76 -438
rect 30 -472 42 -438
rect -88 -478 -30 -472
rect 30 -478 88 -472
<< pwell >>
rect -285 -610 285 610
<< nmos >>
rect -89 -400 -29 400
rect 29 -400 89 400
<< ndiff >>
rect -147 388 -89 400
rect -147 -388 -135 388
rect -101 -388 -89 388
rect -147 -400 -89 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 89 388 147 400
rect 89 -388 101 388
rect 135 -388 147 388
rect 89 -400 147 -388
<< ndiffc >>
rect -135 -388 -101 388
rect -17 -388 17 388
rect 101 -388 135 388
<< psubdiff >>
rect -249 540 -153 574
rect 153 540 249 574
rect -249 478 -215 540
rect 215 478 249 540
rect -249 -540 -215 -478
rect 215 -540 249 -478
rect -249 -574 -153 -540
rect 153 -574 249 -540
<< psubdiffcont >>
rect -153 540 153 574
rect -249 -478 -215 478
rect 215 -478 249 478
rect -153 -574 153 -540
<< poly >>
rect -92 472 -26 488
rect -92 438 -76 472
rect -42 438 -26 472
rect -92 422 -26 438
rect 26 472 92 488
rect 26 438 42 472
rect 76 438 92 472
rect 26 422 92 438
rect -89 400 -29 422
rect 29 400 89 422
rect -89 -422 -29 -400
rect 29 -422 89 -400
rect -92 -438 -26 -422
rect -92 -472 -76 -438
rect -42 -472 -26 -438
rect -92 -488 -26 -472
rect 26 -438 92 -422
rect 26 -472 42 -438
rect 76 -472 92 -438
rect 26 -488 92 -472
<< polycont >>
rect -76 438 -42 472
rect 42 438 76 472
rect -76 -472 -42 -438
rect 42 -472 76 -438
<< locali >>
rect -249 540 -153 574
rect 153 540 249 574
rect -249 478 -215 540
rect 215 478 249 540
rect -92 438 -76 472
rect -42 438 -26 472
rect 26 438 42 472
rect 76 438 92 472
rect -135 388 -101 404
rect -135 -404 -101 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 101 388 135 404
rect 101 -404 135 -388
rect -92 -472 -76 -438
rect -42 -472 -26 -438
rect 26 -472 42 -438
rect 76 -472 92 -438
rect -249 -540 -215 -478
rect 215 -540 249 -478
rect -249 -574 -153 -540
rect 153 -574 249 -540
<< viali >>
rect -76 438 -42 472
rect 42 438 76 472
rect -135 -388 -101 388
rect -17 -388 17 388
rect 101 -388 135 388
rect -76 -472 -42 -438
rect 42 -472 76 -438
<< metal1 >>
rect -88 472 -30 478
rect -88 438 -76 472
rect -42 438 -30 472
rect -88 432 -30 438
rect 30 472 88 478
rect 30 438 42 472
rect 76 438 88 472
rect 30 432 88 438
rect -141 388 -95 400
rect -141 -388 -135 388
rect -101 -388 -95 388
rect -141 -400 -95 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 95 388 141 400
rect 95 -388 101 388
rect 135 -388 141 388
rect 95 -400 141 -388
rect -88 -438 -30 -432
rect -88 -472 -76 -438
rect -42 -472 -30 -438
rect -88 -478 -30 -472
rect 30 -438 88 -432
rect 30 -472 42 -438
rect 76 -472 88 -438
rect 30 -478 88 -472
<< properties >>
string FIXED_BBOX -232 -557 232 557
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.0 l 0.3 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
