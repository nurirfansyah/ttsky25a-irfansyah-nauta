magic
tech sky130A
timestamp 1757964080
<< metal1 >>
rect 5630 4170 5795 4195
rect 5630 4080 5650 4170
rect 5770 4080 5795 4170
rect 5630 4040 5795 4080
rect 6905 4115 7005 4135
rect 6905 4050 6920 4115
rect 6980 4050 7005 4115
rect 6905 4035 7005 4050
rect 7060 4125 7160 4140
rect 7060 4060 7085 4125
rect 7145 4060 7160 4125
rect 7060 4040 7160 4060
rect 7865 4125 7965 4140
rect 7865 4050 7875 4125
rect 7940 4050 7965 4125
rect 7865 4040 7965 4050
rect 8040 4130 8140 4145
rect 8040 4060 8050 4130
rect 8120 4060 8140 4130
rect 8040 4045 8140 4060
rect 4910 3915 8620 3985
rect 4910 3650 5130 3915
rect 5365 3650 8620 3915
rect 4910 3615 8620 3650
rect 5285 2885 6210 3615
rect 7180 2450 8450 3615
rect 8040 2345 8150 2360
rect 8040 2275 8055 2345
rect 8130 2275 8150 2345
rect 8040 2255 8150 2275
rect 7055 2180 7155 2205
rect 7055 2095 7070 2180
rect 7130 2095 7155 2180
rect 7055 2075 7155 2095
rect 6270 1790 6455 1830
rect 4690 1630 4855 1770
rect 5680 1755 5855 1775
rect 5150 1655 5535 1755
rect 5595 1725 6035 1755
rect 5595 1655 5710 1725
rect 5680 1610 5710 1655
rect 5800 1655 6035 1725
rect 6270 1655 6300 1790
rect 6390 1655 6455 1790
rect 7500 1765 7610 1785
rect 5800 1610 5855 1655
rect 5680 1545 5855 1610
rect 6270 1595 6455 1655
rect 6740 1675 7150 1755
rect 6740 1495 6830 1675
rect 7500 1670 7520 1765
rect 7585 1670 7610 1765
rect 8470 1755 8580 1770
rect 7685 1715 8135 1730
rect 7500 1630 7610 1670
rect 7680 1660 8135 1715
rect 8470 1660 8490 1755
rect 8555 1660 8580 1755
rect 6725 1450 6850 1495
rect 6725 1375 6750 1450
rect 6815 1375 6850 1450
rect 6725 1330 6850 1375
rect 6905 1470 7015 1495
rect 6905 1370 6915 1470
rect 6990 1445 7015 1470
rect 7680 1445 7800 1660
rect 8470 1615 8580 1660
rect 6990 1370 7150 1445
rect 6905 1365 7150 1370
rect 7680 1370 7695 1445
rect 7755 1370 7800 1445
rect 6905 1335 7015 1365
rect 7680 1335 7800 1370
rect 7865 1300 8165 1310
rect 7865 1230 7880 1300
rect 7955 1230 8165 1300
rect 7865 1215 8165 1230
rect 5285 655 6230 920
rect 7175 655 8415 1110
rect 4920 100 8615 655
rect 5285 -145 6230 100
rect 7175 -225 8415 100
rect 7845 -390 7970 -360
rect 7845 -455 7850 -390
rect 7950 -455 8140 -390
rect 7845 -470 8140 -455
rect 7850 -480 7955 -470
rect 6770 -575 6900 -545
rect 6770 -640 6800 -575
rect 6880 -640 6900 -575
rect 7010 -550 7120 -525
rect 7010 -615 7030 -550
rect 7090 -615 7120 -550
rect 7010 -630 7120 -615
rect 7680 -570 7780 -550
rect 6770 -675 6900 -640
rect 7680 -640 7700 -570
rect 7760 -640 7780 -570
rect 7680 -665 7780 -640
rect 5665 -815 5850 -765
rect 4725 -1015 4890 -875
rect 5665 -900 5695 -815
rect 5170 -950 5695 -900
rect 5785 -900 5850 -815
rect 6340 -835 6515 -790
rect 5785 -950 6020 -900
rect 5170 -1000 6020 -950
rect 6340 -950 6385 -835
rect 6475 -950 6515 -835
rect 6795 -825 6890 -675
rect 7530 -815 7625 -795
rect 6795 -935 7140 -825
rect 7530 -920 7550 -815
rect 7605 -920 7625 -815
rect 7695 -815 7765 -665
rect 8470 -815 8565 -785
rect 7695 -885 8125 -815
rect 7695 -890 7765 -885
rect 7530 -940 7625 -920
rect 8470 -895 8485 -815
rect 8545 -895 8565 -815
rect 8470 -930 8565 -895
rect 6340 -1020 6515 -950
rect 7025 -1280 7145 -1260
rect 7025 -1375 7040 -1280
rect 7130 -1375 7145 -1280
rect 7025 -1400 7145 -1375
rect 8025 -1405 8150 -1380
rect 8025 -1495 8045 -1405
rect 8125 -1495 8150 -1405
rect 8025 -1515 8150 -1495
rect 5280 -2870 6200 -2085
rect 7205 -2870 8450 -1620
rect 4910 -2900 8615 -2870
rect 4910 -3165 5140 -2900
rect 5375 -3165 8615 -2900
rect 4910 -3215 8615 -3165
rect 6720 -3300 6855 -3265
rect 5615 -3405 5840 -3380
rect 6720 -3385 6730 -3300
rect 6825 -3385 6855 -3300
rect 7035 -3285 7135 -3270
rect 7035 -3365 7045 -3285
rect 7120 -3365 7135 -3285
rect 7845 -3280 7945 -3260
rect 7845 -3350 7855 -3280
rect 7920 -3350 7945 -3280
rect 7845 -3360 7945 -3350
rect 7995 -3285 8095 -3270
rect 7995 -3355 8010 -3285
rect 8070 -3355 8095 -3285
rect 7035 -3370 7135 -3365
rect 7995 -3370 8095 -3355
rect 6720 -3400 6855 -3385
rect 5615 -3490 5660 -3405
rect 5805 -3490 5840 -3405
rect 5615 -3520 5840 -3490
<< via1 >>
rect 5650 4080 5770 4170
rect 6920 4050 6980 4115
rect 7085 4060 7145 4125
rect 7875 4050 7940 4125
rect 8050 4060 8120 4130
rect 5130 3650 5365 3915
rect 8055 2275 8130 2345
rect 7070 2095 7130 2180
rect 5710 1610 5800 1725
rect 6300 1655 6390 1790
rect 7520 1670 7585 1765
rect 8490 1660 8555 1755
rect 6750 1375 6815 1450
rect 6915 1370 6990 1470
rect 7695 1370 7755 1445
rect 7880 1230 7955 1300
rect 7850 -455 7950 -390
rect 6800 -640 6880 -575
rect 7030 -615 7090 -550
rect 7700 -640 7760 -570
rect 5695 -950 5785 -815
rect 6385 -950 6475 -835
rect 7550 -920 7605 -815
rect 8485 -895 8545 -815
rect 7040 -1375 7130 -1280
rect 8045 -1495 8125 -1405
rect 5140 -3165 5375 -2900
rect 6730 -3385 6825 -3300
rect 7045 -3365 7120 -3285
rect 7855 -3350 7920 -3280
rect 8010 -3355 8070 -3285
rect 5660 -3490 5805 -3405
<< metal2 >>
rect 5630 4170 5795 4195
rect 5630 4080 5650 4170
rect 5770 4080 5795 4170
rect 5115 3915 5385 3935
rect 5115 3650 5130 3915
rect 5365 3650 5385 3915
rect 5115 -2880 5385 3650
rect 5630 2050 5795 4080
rect 6905 4115 7005 4135
rect 6905 4050 6920 4115
rect 6980 4050 7005 4115
rect 6905 4035 7005 4050
rect 6515 2050 6675 2055
rect 5630 1950 6680 2050
rect 5685 1880 6680 1950
rect 5685 1775 5835 1880
rect 6270 1790 6455 1830
rect 5680 1725 5855 1775
rect 5680 1640 5710 1725
rect 5670 1610 5710 1640
rect 5800 1610 5855 1725
rect 5670 1545 5855 1610
rect 6270 1655 6300 1790
rect 6390 1655 6455 1790
rect 6270 1595 6455 1655
rect 5670 1445 5830 1545
rect 5670 1375 5710 1445
rect 5785 1375 5830 1445
rect 5670 1330 5830 1375
rect 6300 915 6435 1595
rect 6300 825 6315 915
rect 6405 825 6435 915
rect 6300 565 6435 825
rect 5700 540 6435 565
rect 5690 375 6435 540
rect 5690 -540 5825 375
rect 6300 370 6435 375
rect 6515 -5 6675 1880
rect 6920 1495 7005 4035
rect 7060 4125 7160 4140
rect 7060 4060 7085 4125
rect 7145 4060 7160 4125
rect 7060 4040 7160 4060
rect 7865 4125 7970 4140
rect 7865 4050 7875 4125
rect 7940 4050 7970 4125
rect 7060 2205 7130 4040
rect 7055 2180 7155 2205
rect 7055 2095 7070 2180
rect 7130 2095 7155 2180
rect 7055 2075 7155 2095
rect 7500 1765 7610 1785
rect 7500 1670 7520 1765
rect 7585 1670 7610 1765
rect 7500 1630 7610 1670
rect 6725 1450 6850 1495
rect 6725 1375 6750 1450
rect 6815 1375 6850 1450
rect 6725 1330 6850 1375
rect 6905 1470 7015 1495
rect 6905 1370 6915 1470
rect 6990 1370 7015 1470
rect 6905 1335 7015 1370
rect 7515 925 7600 1630
rect 7685 1445 7795 1505
rect 7685 1370 7695 1445
rect 7755 1370 7795 1445
rect 7685 1345 7795 1370
rect 7865 1300 7970 4050
rect 8040 4130 8145 4150
rect 8040 4060 8050 4130
rect 8120 4060 8145 4130
rect 8040 2360 8145 4060
rect 8040 2345 8150 2360
rect 8040 2275 8055 2345
rect 8130 2275 8150 2345
rect 8040 2255 8150 2275
rect 8470 1755 8580 1770
rect 8470 1660 8490 1755
rect 8555 1660 8580 1755
rect 8470 1615 8580 1660
rect 7865 1230 7880 1300
rect 7955 1230 7970 1300
rect 7865 1215 7970 1230
rect 8480 925 8565 1615
rect 6810 910 8565 925
rect 6810 820 6840 910
rect 6930 885 8565 910
rect 6930 820 8560 885
rect 6810 815 8560 820
rect 6515 -110 8615 -5
rect 5690 -575 5835 -540
rect 5690 -640 5715 -575
rect 5795 -640 5835 -575
rect 5690 -665 5835 -640
rect 5690 -765 5825 -665
rect 5665 -775 5850 -765
rect 5615 -815 5850 -775
rect 6515 -790 6675 -110
rect 7010 -550 7120 -525
rect 6760 -575 6900 -550
rect 6760 -640 6800 -575
rect 6880 -640 6900 -575
rect 6760 -675 6900 -640
rect 7010 -615 7030 -550
rect 7090 -615 7120 -550
rect 7010 -630 7120 -615
rect 5615 -950 5695 -815
rect 5785 -950 5850 -815
rect 5615 -1000 5850 -950
rect 6340 -835 6675 -790
rect 6340 -950 6385 -835
rect 6475 -950 6675 -835
rect 5115 -2900 5405 -2880
rect 5115 -3165 5140 -2900
rect 5375 -3165 5405 -2900
rect 5115 -3205 5405 -3165
rect 5615 -3405 5840 -1000
rect 6340 -1015 6675 -950
rect 6340 -1020 6515 -1015
rect 7010 -1090 7100 -630
rect 7550 -795 7625 -110
rect 7845 -390 7970 -365
rect 7845 -455 7850 -390
rect 7950 -455 7970 -390
rect 7845 -480 7970 -455
rect 7680 -570 7780 -550
rect 7680 -640 7700 -570
rect 7760 -640 7780 -570
rect 7680 -665 7780 -640
rect 7530 -815 7625 -795
rect 7530 -920 7550 -815
rect 7605 -920 7625 -815
rect 7530 -940 7625 -920
rect 6735 -1165 7100 -1090
rect 6735 -3265 6825 -1165
rect 7025 -1280 7145 -1260
rect 7025 -1375 7040 -1280
rect 7130 -1375 7145 -1280
rect 6720 -3300 6855 -3265
rect 6720 -3385 6730 -3300
rect 6825 -3385 6855 -3300
rect 6720 -3400 6855 -3385
rect 7025 -3285 7145 -1375
rect 7860 -3260 7940 -480
rect 8540 -785 8615 -110
rect 8470 -815 8615 -785
rect 8470 -895 8485 -815
rect 8545 -855 8615 -815
rect 8545 -895 8565 -855
rect 8470 -930 8565 -895
rect 8025 -1405 8150 -1380
rect 8025 -1420 8045 -1405
rect 8020 -1495 8045 -1420
rect 8125 -1495 8150 -1405
rect 8020 -1515 8150 -1495
rect 7025 -3365 7045 -3285
rect 7120 -3365 7145 -3285
rect 7845 -3280 7945 -3260
rect 8020 -3270 8090 -1515
rect 7845 -3350 7855 -3280
rect 7920 -3350 7945 -3280
rect 7845 -3360 7945 -3350
rect 7995 -3285 8095 -3270
rect 7995 -3355 8010 -3285
rect 8070 -3355 8095 -3285
rect 7025 -3390 7145 -3365
rect 7995 -3370 8095 -3355
rect 5615 -3490 5660 -3405
rect 5805 -3490 5840 -3405
rect 5615 -3520 5840 -3490
<< via2 >>
rect 5710 1375 5785 1445
rect 6315 825 6405 915
rect 6750 1375 6815 1450
rect 7695 1370 7755 1445
rect 6840 820 6930 910
rect 5715 -640 5795 -575
rect 6800 -640 6880 -575
rect 7700 -640 7760 -570
<< metal3 >>
rect 5665 1450 7780 1475
rect 5665 1445 6750 1450
rect 5665 1375 5710 1445
rect 5785 1375 6750 1445
rect 6815 1445 7780 1450
rect 6815 1375 7695 1445
rect 5665 1370 7695 1375
rect 7755 1370 7780 1445
rect 5665 1340 7780 1370
rect 6295 915 6950 955
rect 6295 825 6315 915
rect 6405 910 6950 915
rect 6405 825 6840 910
rect 6295 820 6840 825
rect 6930 820 6950 910
rect 6295 795 6950 820
rect 5695 -565 5835 -540
rect 7680 -565 7780 -550
rect 5695 -570 7780 -565
rect 5695 -575 7700 -570
rect 5695 -640 5715 -575
rect 5795 -640 6800 -575
rect 6880 -640 7700 -575
rect 7760 -640 7780 -570
rect 5695 -660 7780 -640
rect 5695 -665 5835 -660
rect 7680 -665 7780 -660
use ff_inv  x1
timestamp 1757958233
transform 1 0 3685 0 1 1755
box 1155 -1195 1565 1920
use ff_inv  x2
timestamp 1757958233
transform 1 0 3705 0 -1 -1000
box 1155 -1195 1565 1920
use sc_inv  x3
timestamp 1757958533
transform 1 0 4730 0 1 2085
box 550 -1275 875 885
use sc_inv  x4
timestamp 1757958533
transform 1 0 4735 0 -1 -1330
box 550 -1275 875 885
use cc_inv_4  x5
timestamp 1757958378
transform 1 0 5595 0 1 1940
box 385 -1095 740 975
use cc_inv_4  x6
timestamp 1757958378
transform 1 0 5610 0 -1 -1185
box 385 -1095 740 975
use cc_inv_dt05  x7
timestamp 1757958777
transform 1 0 6595 0 1 2215
box 490 -1195 930 260
use cc_inv_dt05  x8
timestamp 1757958777
transform 1 0 6605 0 -1 -1395
box 490 -1195 930 260
use cc_inv_dt05_long  x11
timestamp 1757958958
transform 1 0 7575 0 1 2095
box 475 -1090 900 450
use cc_inv_dt05_long  x12
timestamp 1757958958
transform 1 0 7575 0 -1 -1260
box 475 -1090 900 450
<< labels >>
flabel metal1 5035 3840 5135 3940 0 FreeSans 128 0 0 0 vdd
port 0 nsew
flabel metal1 5090 305 5190 405 0 FreeSans 128 0 0 0 gnd
port 13 nsew
flabel metal1 4700 1660 4800 1760 0 FreeSans 128 0 0 0 in_p
port 2 nsew
flabel metal1 4725 -1000 4825 -900 0 FreeSans 128 0 0 0 in_n
port 4 nsew
flabel metal1 5650 4045 5750 4145 0 FreeSans 128 0 0 0 out_n
port 1 nsew
flabel metal1 5625 -3485 5725 -3385 0 FreeSans 128 0 0 0 out_p
port 3 nsew
flabel metal1 7060 4040 7160 4140 0 FreeSans 128 0 0 0 sw_p_A1
port 5 nsew
flabel metal1 6905 4035 7005 4135 0 FreeSans 128 0 0 0 sw_n_A1
port 9 nsew
flabel metal1 7865 4040 7965 4140 0 FreeSans 128 0 0 0 sw_n_A05
port 11 nsew
flabel metal1 8040 4045 8140 4145 0 FreeSans 128 0 0 0 sw_p_A05
port 7 nsew
flabel metal1 7035 -3370 7135 -3270 0 FreeSans 128 0 0 0 sw_p_B1
port 6 nsew
flabel metal1 6735 -3375 6835 -3275 0 FreeSans 128 0 0 0 sw_n_B1
port 10 nsew
flabel metal1 7995 -3370 8095 -3270 0 FreeSans 128 0 0 0 sw_p_B05
port 8 nsew
flabel metal1 7845 -3360 7945 -3260 0 FreeSans 128 0 0 0 sw_n_B05
port 12 nsew
<< end >>
