** sch_path: /home/irfansyah/design/ttsky25a-irfansyah-nauta/xsch/tt_um_nurirfansyah_nauta.sch
**.subckt tt_um_nurirfansyah_nauta clk ena rst_n ua[3] ua[4] ua[5] ua[6] ua[7] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5]
*+ ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3]
*+ uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] uio_out[0] uio_out[1]
*+ uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] ua[2] ua[1] ui_in[0] uo_out[0] ua[0] VGND VPWR
*.ipin clk
*.ipin ena
*.ipin rst_n
*.opin ua[3]
*.ipin ua[4]
*.ipin ua[5]
*.ipin ua[6]
*.ipin ua[7]
*.ipin ui_in[1]
*.ipin ui_in[2]
*.ipin ui_in[3]
*.ipin ui_in[4]
*.ipin ui_in[5]
*.ipin ui_in[6]
*.ipin ui_in[7]
*.ipin uio_in[0]
*.ipin uio_in[1]
*.ipin uio_in[2]
*.ipin uio_in[3]
*.ipin uio_in[4]
*.ipin uio_in[5]
*.ipin uio_in[6]
*.ipin uio_in[7]
*.opin uio_oe[0]
*.opin uio_oe[1]
*.opin uio_oe[2]
*.opin uio_oe[3]
*.opin uio_oe[4]
*.opin uio_oe[5]
*.opin uio_oe[6]
*.opin uio_oe[7]
*.opin uo_out[1]
*.opin uo_out[2]
*.opin uo_out[3]
*.opin uo_out[4]
*.opin uo_out[5]
*.opin uo_out[6]
*.opin uo_out[7]
*.iopin uio_out[0]
*.iopin uio_out[1]
*.iopin uio_out[2]
*.iopin uio_out[3]
*.iopin uio_out[4]
*.iopin uio_out[5]
*.iopin uio_out[6]
*.iopin uio_out[7]
*.opin ua[2]
*.ipin ua[1]
*.ipin ui_in[0]
*.opin uo_out[0]
*.ipin ua[0]
*.iopin VGND
*.iopin VPWR
* noconn clk
* noconn ena
* noconn rst_n
* noconn ua[6]
* noconn uio_in[0]
* noconn uio_in[1]
* noconn uio_in[2]
* noconn uio_in[3]
* noconn uio_in[4]
* noconn uio_in[5]
* noconn uio_in[6]
* noconn uio_in[7]
* noconn ua[5]
* noconn ua[4]
* noconn ua[7]
* noconn uio_oe[0]
* noconn uio_oe[1]
* noconn uio_oe[2]
* noconn uio_oe[3]
* noconn uio_oe[4]
* noconn uio_oe[5]
* noconn uio_oe[6]
* noconn uio_oe[7]
* noconn uo_out[5]
* noconn uo_out[6]
* noconn uo_out[7]
* noconn uio_out[0]
* noconn uio_out[1]
* noconn uio_out[2]
* noconn uio_out[3]
* noconn uio_out[4]
* noconn uio_out[5]
* noconn uio_out[6]
* noconn uio_out[7]
x1 VPWR ua[2] ua[0] ua[3] ua[1] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] VGND nauta_ota_dtrim2b
* noconn uo_out[0]
* noconn uo_out[1]
* noconn uo_out[2]
* noconn uo_out[3]
* noconn uo_out[4]
**.ends

* expanding   symbol:  nauta_ota_dtrim2b.sym # of pins=14
** sym_path: /home/irfansyah/design/ttsky25a-irfansyah-nauta/xsch/nauta_ota_dtrim2b.sym
** sch_path: /home/irfansyah/design/ttsky25a-irfansyah-nauta/xsch/nauta_ota_dtrim2b.sch
.subckt nauta_ota_dtrim2b vdd out_n in_p out_p in_n sw_p_A1 sw_p_B1 sw_p_A05 sw_p_B05 sw_n_A1 sw_n_B1 sw_n_A05 sw_n_B05 gnd
*.ipin vdd
*.ipin gnd
*.ipin in_n
*.ipin in_p
*.opin out_n
*.opin out_p
*.ipin sw_p_A05
*.ipin sw_n_B1
*.ipin sw_p_A1
*.ipin sw_p_B1
*.ipin sw_p_B05
*.ipin sw_n_A1
*.ipin sw_n_A05
*.ipin sw_n_B05
x1 vdd in_p out_n gnd ff_inv
x2 vdd in_n out_p gnd ff_inv
x3 vdd out_n out_n gnd sc_inv
x4 vdd out_p out_p gnd sc_inv
x5 vdd out_n out_p gnd cc_inv_4
x6 vdd out_p out_n gnd cc_inv_4
x7 vdd out_p out_n sw_p_A1 sw_n_A1 gnd cc_inv_dt05
x8 vdd out_n out_p sw_p_B1 sw_n_B1 gnd cc_inv_dt05
x11 vdd out_p out_n sw_p_A05 sw_n_A05 gnd cc_inv_dt05_long
x12 vdd out_n out_p sw_p_B05 sw_n_B05 gnd cc_inv_dt05_long
.ends


* expanding   symbol:  ff_inv.sym # of pins=4
** sym_path: /home/irfansyah/design/ttsky25a-irfansyah-nauta/xsch/ff_inv.sym
** sch_path: /home/irfansyah/design/ttsky25a-irfansyah-nauta/xsch/ff_inv.sch
.subckt ff_inv vdd in out gnd
*.ipin in
*.ipin vdd
*.ipin gnd
*.opin out
XM1 out in gnd gnd sky130_fd_pr__nfet_01v8 L=0.3 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  sc_inv.sym # of pins=4
** sym_path: /home/irfansyah/design/ttsky25a-irfansyah-nauta/xsch/sc_inv.sym
** sch_path: /home/irfansyah/design/ttsky25a-irfansyah-nauta/xsch/sc_inv.sch
.subckt sc_inv vdd in out gnd
*.ipin in
*.ipin vdd
*.ipin gnd
*.opin out
XM1 out in gnd gnd sky130_fd_pr__nfet_01v8 L=0.3 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  cc_inv_4.sym # of pins=4
** sym_path: /home/irfansyah/design/ttsky25a-irfansyah-nauta/xsch/cc_inv_4.sym
** sch_path: /home/irfansyah/design/ttsky25a-irfansyah-nauta/xsch/cc_inv_4.sch
.subckt cc_inv_4 vdd in out gnd
*.ipin in
*.ipin vdd
*.ipin gnd
*.opin out
XM1 out in gnd gnd sky130_fd_pr__nfet_01v8 L=0.3 W=3.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=7.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  cc_inv_dt05.sym # of pins=6
** sym_path: /home/irfansyah/design/ttsky25a-irfansyah-nauta/xsch/cc_inv_dt05.sym
** sch_path: /home/irfansyah/design/ttsky25a-irfansyah-nauta/xsch/cc_inv_dt05.sch
.subckt cc_inv_dt05 vdd out in sw_p sw_n gnd
*.ipin in
*.ipin vdd
*.ipin gnd
*.opin out
*.ipin sw_n
*.ipin sw_p
XM1 out in net1 gnd sky130_fd_pr__nfet_01v8 L=0.3 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in net2 vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 sw_p vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 sw_n gnd gnd sky130_fd_pr__nfet_01v8 L=0.3 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  cc_inv_dt05_long.sym # of pins=6
** sym_path: /home/irfansyah/design/ttsky25a-irfansyah-nauta/xsch/cc_inv_dt05_long.sym
** sch_path: /home/irfansyah/design/ttsky25a-irfansyah-nauta/xsch/cc_inv_dt05_long.sch
.subckt cc_inv_dt05_long vdd out in sw_p sw_n gnd
*.ipin in
*.ipin vdd
*.ipin gnd
*.opin out
*.ipin sw_n
*.ipin sw_p
XM1 out in net1 gnd sky130_fd_pr__nfet_01v8 L=0.4 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in net2 vdd sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 sw_p vdd vdd sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 sw_n gnd gnd sky130_fd_pr__nfet_01v8 L=0.4 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
