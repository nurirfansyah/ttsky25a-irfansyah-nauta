magic
tech sky130A
magscale 1 2
timestamp 1757958233
<< locali >>
rect 2460 3620 2930 3640
rect 2460 3570 2490 3620
rect 2900 3570 2930 3620
rect 2460 3550 2930 3570
rect 2470 -2140 2920 -2130
rect 2470 -2190 2490 -2140
rect 2900 -2190 2920 -2140
rect 2470 -2200 2920 -2190
<< viali >>
rect 2490 3570 2900 3620
rect 2490 -2190 2900 -2140
<< metal1 >>
rect 2460 3620 2930 3840
rect 2460 3570 2490 3620
rect 2900 3570 2930 3620
rect 2460 3550 2930 3570
rect 2550 3340 2620 3550
rect 2660 3470 2740 3520
rect 2310 -40 2510 0
rect 2660 -40 2730 170
rect 2310 -130 2730 -40
rect 2310 -200 2510 -130
rect 2660 -270 2730 -130
rect 2650 -350 2730 -270
rect 2770 -40 2810 290
rect 2930 -40 3130 0
rect 2770 -130 3130 -40
rect 2770 -470 2810 -130
rect 2930 -200 3130 -130
rect 2572 -2130 2614 -1894
rect 2660 -2086 2728 -2018
rect 2470 -2140 2930 -2130
rect 2470 -2190 2490 -2140
rect 2900 -2190 2930 -2140
rect 2470 -2390 2930 -2190
use sky130_fd_pr__nfet_01v8_RMGWKL  XM1
timestamp 1757952087
transform 1 0 2696 0 1 -1180
box -226 -1010 226 1010
use sky130_fd_pr__pfet_01v8_XP7VY6  XM2
timestamp 1757952087
transform 1 0 2696 0 1 1829
box -226 -1819 226 1819
<< labels >>
flabel metal1 2460 3640 2660 3840 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 2470 -2390 2670 -2190 0 FreeSans 256 0 0 0 gnd
port 3 nsew
flabel metal1 2310 -200 2510 0 0 FreeSans 256 0 0 0 in
port 1 nsew
flabel metal1 2930 -200 3130 0 0 FreeSans 256 0 0 0 out
port 2 nsew
<< end >>
