VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_sky25a_nurirfansyah_nauta
  CLASS BLOCK ;
  FOREIGN tt_um_sky25a_nurirfansyah_nauta ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.070000 ;
    ANTENNADIFFAREA 14.615999 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.070000 ;
    ANTENNADIFFAREA 14.615999 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.400000 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.400000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.150000 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.150000 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.200000 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.200000 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT -0.600 80.250 0.000 92.000 ;
        RECT -0.300 24.400 0.000 35.950 ;
      LAYER met2 ;
        RECT -0.600 80.250 0.000 92.000 ;
        RECT -0.300 24.400 0.000 35.950 ;
      LAYER met3 ;
        RECT -0.600 80.250 0.000 92.000 ;
        RECT -0.300 24.400 0.000 35.950 ;
      LAYER met4 ;
        RECT -0.600 80.250 0.000 92.000 ;
        RECT -0.300 24.400 0.000 35.950 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 100.090 72.450 102.740 79.400 ;
        RECT 110.190 72.300 112.590 78.950 ;
        RECT 122.430 73.150 124.690 82.940 ;
        RECT 129.330 73.150 131.590 83.340 ;
        RECT 133.080 72.600 135.340 90.790 ;
      LAYER pwell ;
        RECT 100.290 68.910 102.650 71.510 ;
        RECT 110.280 69.150 112.540 71.750 ;
        RECT 100.300 66.150 102.660 68.750 ;
        RECT 110.290 68.700 112.540 69.150 ;
        RECT 110.230 68.650 112.540 68.700 ;
        RECT 110.230 66.100 112.490 68.650 ;
        RECT 122.430 64.650 124.690 70.550 ;
        RECT 129.330 64.400 131.590 70.500 ;
        RECT 133.080 61.600 135.340 71.700 ;
        RECT 100.300 49.600 102.660 52.200 ;
        RECT 110.130 49.550 112.390 52.100 ;
        RECT 110.130 49.500 112.440 49.550 ;
        RECT 100.290 46.840 102.650 49.440 ;
        RECT 110.190 49.050 112.440 49.500 ;
        RECT 110.180 46.450 112.440 49.050 ;
        RECT 122.280 47.000 124.540 52.900 ;
        RECT 129.280 47.050 131.540 53.150 ;
      LAYER nwell ;
        RECT 100.090 38.950 102.740 45.900 ;
        RECT 110.090 39.250 112.490 45.900 ;
      LAYER pwell ;
        RECT 132.880 45.850 135.140 55.950 ;
      LAYER nwell ;
        RECT 122.280 34.610 124.540 44.400 ;
        RECT 129.280 34.210 131.540 44.400 ;
        RECT 132.880 26.760 135.140 44.950 ;
      LAYER li1 ;
        RECT 133.040 90.300 135.390 90.750 ;
        RECT 122.440 82.600 124.690 83.150 ;
        RECT 129.290 82.950 131.640 83.450 ;
        RECT 122.610 82.590 124.510 82.600 ;
        RECT 100.090 79.000 102.740 79.450 ;
        RECT 100.420 76.520 100.590 79.000 ;
        RECT 101.220 78.500 101.620 78.670 ;
        RECT 100.990 77.245 101.160 78.285 ;
        RECT 101.680 77.245 101.850 78.285 ;
        RECT 101.220 76.860 101.620 77.030 ;
        RECT 102.250 76.520 102.420 79.000 ;
        RECT 110.190 78.500 112.590 78.900 ;
        RECT 100.420 76.350 102.420 76.520 ;
        RECT 110.460 78.440 112.360 78.500 ;
        RECT 100.890 75.600 101.940 76.350 ;
        RECT 110.460 75.950 110.630 78.440 ;
        RECT 111.245 77.930 111.575 78.100 ;
        RECT 111.030 76.675 111.200 77.715 ;
        RECT 111.620 76.675 111.790 77.715 ;
        RECT 111.245 76.290 111.575 76.460 ;
        RECT 112.190 75.950 112.360 78.440 ;
        RECT 110.460 75.780 112.360 75.950 ;
        RECT 100.440 75.430 102.440 75.600 ;
        RECT 100.440 72.940 100.610 75.430 ;
        RECT 101.240 74.920 101.640 75.090 ;
        RECT 101.010 73.665 101.180 74.705 ;
        RECT 101.700 73.665 101.870 74.705 ;
        RECT 101.240 73.280 101.640 73.450 ;
        RECT 102.270 72.940 102.440 75.430 ;
        RECT 110.640 75.360 112.190 75.780 ;
        RECT 100.440 72.770 102.440 72.940 ;
        RECT 110.460 75.190 112.360 75.360 ;
        RECT 110.460 72.700 110.630 75.190 ;
        RECT 111.245 74.680 111.575 74.850 ;
        RECT 111.030 73.425 111.200 74.465 ;
        RECT 111.620 73.425 111.790 74.465 ;
        RECT 111.245 73.040 111.575 73.210 ;
        RECT 112.190 72.700 112.360 75.190 ;
        RECT 122.610 73.500 122.780 82.590 ;
        RECT 123.395 82.080 123.725 82.250 ;
        RECT 123.180 74.225 123.350 81.865 ;
        RECT 123.770 74.225 123.940 81.865 ;
        RECT 123.395 73.840 123.725 74.010 ;
        RECT 124.340 73.500 124.510 82.590 ;
        RECT 122.610 73.330 124.510 73.500 ;
        RECT 129.510 73.500 129.680 82.950 ;
        RECT 130.295 82.480 130.625 82.650 ;
        RECT 130.080 74.225 130.250 82.265 ;
        RECT 130.670 74.225 130.840 82.265 ;
        RECT 130.295 73.840 130.625 74.010 ;
        RECT 131.240 73.500 131.410 82.950 ;
        RECT 129.510 73.330 131.410 73.500 ;
        RECT 133.260 72.950 133.430 90.300 ;
        RECT 134.045 89.930 134.375 90.100 ;
        RECT 133.830 73.675 134.000 89.715 ;
        RECT 134.420 73.675 134.590 89.715 ;
        RECT 134.045 73.290 134.375 73.460 ;
        RECT 134.990 72.950 135.160 90.300 ;
        RECT 133.260 72.780 135.160 72.950 ;
        RECT 110.460 72.530 112.360 72.700 ;
        RECT 110.460 71.400 112.360 71.570 ;
        RECT 100.470 71.160 102.470 71.330 ;
        RECT 100.470 69.260 100.640 71.160 ;
        RECT 101.270 70.650 101.670 70.820 ;
        RECT 101.040 69.940 101.210 70.480 ;
        RECT 101.730 69.940 101.900 70.480 ;
        RECT 101.270 69.600 101.670 69.770 ;
        RECT 102.300 69.260 102.470 71.160 ;
        RECT 110.460 69.500 110.630 71.400 ;
        RECT 111.245 70.890 111.575 71.060 ;
        RECT 111.030 70.180 111.200 70.720 ;
        RECT 111.620 70.180 111.790 70.720 ;
        RECT 111.245 69.840 111.575 70.010 ;
        RECT 112.190 69.500 112.360 71.400 ;
        RECT 133.260 71.350 135.160 71.520 ;
        RECT 110.460 69.330 112.360 69.500 ;
        RECT 122.610 70.200 124.510 70.370 ;
        RECT 100.470 69.090 102.470 69.260 ;
        RECT 101.090 68.570 101.790 69.090 ;
        RECT 100.480 68.400 102.480 68.570 ;
        RECT 100.480 66.500 100.650 68.400 ;
        RECT 101.280 67.890 101.680 68.060 ;
        RECT 101.050 67.180 101.220 67.720 ;
        RECT 101.740 67.180 101.910 67.720 ;
        RECT 101.280 66.840 101.680 67.010 ;
        RECT 102.310 66.500 102.480 68.400 ;
        RECT 110.410 68.350 112.310 68.520 ;
        RECT 100.290 65.900 102.640 66.500 ;
        RECT 110.410 66.450 110.580 68.350 ;
        RECT 111.195 67.840 111.525 68.010 ;
        RECT 110.980 67.130 111.150 67.670 ;
        RECT 111.570 67.130 111.740 67.670 ;
        RECT 111.195 66.790 111.525 66.960 ;
        RECT 112.140 66.450 112.310 68.350 ;
        RECT 110.240 65.950 112.640 66.450 ;
        RECT 122.610 65.000 122.780 70.200 ;
        RECT 123.395 69.690 123.725 69.860 ;
        RECT 123.180 65.680 123.350 69.520 ;
        RECT 123.770 65.680 123.940 69.520 ;
        RECT 123.395 65.340 123.725 65.510 ;
        RECT 124.340 65.000 124.510 70.200 ;
        RECT 129.510 70.150 131.410 70.320 ;
        RECT 122.390 64.400 124.690 65.000 ;
        RECT 129.510 64.750 129.680 70.150 ;
        RECT 130.295 69.640 130.625 69.810 ;
        RECT 130.080 65.430 130.250 69.470 ;
        RECT 130.670 65.430 130.840 69.470 ;
        RECT 130.295 65.090 130.625 65.260 ;
        RECT 131.240 64.750 131.410 70.150 ;
        RECT 129.290 64.150 131.590 64.750 ;
        RECT 133.260 61.950 133.430 71.350 ;
        RECT 134.045 70.840 134.375 71.010 ;
        RECT 133.830 62.630 134.000 70.670 ;
        RECT 134.420 62.630 134.590 70.670 ;
        RECT 134.045 62.290 134.375 62.460 ;
        RECT 134.990 61.950 135.160 71.350 ;
        RECT 133.260 61.900 135.160 61.950 ;
        RECT 133.090 61.550 135.340 61.900 ;
        RECT 132.890 55.650 135.140 56.000 ;
        RECT 133.060 55.600 134.960 55.650 ;
        RECT 122.240 52.550 124.540 53.150 ;
        RECT 129.240 52.800 131.540 53.400 ;
        RECT 100.290 51.850 102.640 52.450 ;
        RECT 100.480 49.950 100.650 51.850 ;
        RECT 101.280 51.340 101.680 51.510 ;
        RECT 101.050 50.630 101.220 51.170 ;
        RECT 101.740 50.630 101.910 51.170 ;
        RECT 101.280 50.290 101.680 50.460 ;
        RECT 102.310 49.950 102.480 51.850 ;
        RECT 110.140 51.750 112.540 52.250 ;
        RECT 100.480 49.780 102.480 49.950 ;
        RECT 110.310 49.850 110.480 51.750 ;
        RECT 111.095 51.240 111.425 51.410 ;
        RECT 110.880 50.530 111.050 51.070 ;
        RECT 111.470 50.530 111.640 51.070 ;
        RECT 111.095 50.190 111.425 50.360 ;
        RECT 112.040 49.850 112.210 51.750 ;
        RECT 101.090 49.260 101.790 49.780 ;
        RECT 110.310 49.680 112.210 49.850 ;
        RECT 100.470 49.090 102.470 49.260 ;
        RECT 100.470 47.190 100.640 49.090 ;
        RECT 101.270 48.580 101.670 48.750 ;
        RECT 101.040 47.870 101.210 48.410 ;
        RECT 101.730 47.870 101.900 48.410 ;
        RECT 101.270 47.530 101.670 47.700 ;
        RECT 102.300 47.190 102.470 49.090 ;
        RECT 100.470 47.020 102.470 47.190 ;
        RECT 110.360 48.700 112.260 48.870 ;
        RECT 110.360 46.800 110.530 48.700 ;
        RECT 111.145 48.190 111.475 48.360 ;
        RECT 110.930 47.480 111.100 48.020 ;
        RECT 111.520 47.480 111.690 48.020 ;
        RECT 111.145 47.140 111.475 47.310 ;
        RECT 112.090 46.800 112.260 48.700 ;
        RECT 122.460 47.350 122.630 52.550 ;
        RECT 123.245 52.040 123.575 52.210 ;
        RECT 123.030 48.030 123.200 51.870 ;
        RECT 123.620 48.030 123.790 51.870 ;
        RECT 123.245 47.690 123.575 47.860 ;
        RECT 124.190 47.350 124.360 52.550 ;
        RECT 122.460 47.180 124.360 47.350 ;
        RECT 129.460 47.400 129.630 52.800 ;
        RECT 130.245 52.290 130.575 52.460 ;
        RECT 130.030 48.080 130.200 52.120 ;
        RECT 130.620 48.080 130.790 52.120 ;
        RECT 130.245 47.740 130.575 47.910 ;
        RECT 131.190 47.400 131.360 52.800 ;
        RECT 129.460 47.230 131.360 47.400 ;
        RECT 110.360 46.630 112.260 46.800 ;
        RECT 133.060 46.200 133.230 55.600 ;
        RECT 133.845 55.090 134.175 55.260 ;
        RECT 133.630 46.880 133.800 54.920 ;
        RECT 134.220 46.880 134.390 54.920 ;
        RECT 133.845 46.540 134.175 46.710 ;
        RECT 134.790 46.200 134.960 55.600 ;
        RECT 133.060 46.030 134.960 46.200 ;
        RECT 100.440 45.410 102.440 45.580 ;
        RECT 100.440 42.920 100.610 45.410 ;
        RECT 101.240 44.900 101.640 45.070 ;
        RECT 101.010 43.645 101.180 44.685 ;
        RECT 101.700 43.645 101.870 44.685 ;
        RECT 101.240 43.260 101.640 43.430 ;
        RECT 102.270 42.920 102.440 45.410 ;
        RECT 100.440 42.750 102.440 42.920 ;
        RECT 110.360 45.500 112.260 45.670 ;
        RECT 110.360 43.010 110.530 45.500 ;
        RECT 111.145 44.990 111.475 45.160 ;
        RECT 110.930 43.735 111.100 44.775 ;
        RECT 111.520 43.735 111.690 44.775 ;
        RECT 111.145 43.350 111.475 43.520 ;
        RECT 112.090 43.010 112.260 45.500 ;
        RECT 133.060 44.600 134.960 44.770 ;
        RECT 110.360 42.840 112.260 43.010 ;
        RECT 122.460 44.050 124.360 44.220 ;
        RECT 100.890 42.000 101.940 42.750 ;
        RECT 110.540 42.420 112.090 42.840 ;
        RECT 110.360 42.250 112.260 42.420 ;
        RECT 100.420 41.830 102.420 42.000 ;
        RECT 100.420 39.350 100.590 41.830 ;
        RECT 101.220 41.320 101.620 41.490 ;
        RECT 100.990 40.065 101.160 41.105 ;
        RECT 101.680 40.065 101.850 41.105 ;
        RECT 101.220 39.680 101.620 39.850 ;
        RECT 102.250 39.350 102.420 41.830 ;
        RECT 110.360 39.760 110.530 42.250 ;
        RECT 111.145 41.740 111.475 41.910 ;
        RECT 110.930 40.485 111.100 41.525 ;
        RECT 111.520 40.485 111.690 41.525 ;
        RECT 111.145 40.100 111.475 40.270 ;
        RECT 112.090 39.760 112.260 42.250 ;
        RECT 110.360 39.700 112.260 39.760 ;
        RECT 100.090 38.900 102.740 39.350 ;
        RECT 110.090 39.300 112.490 39.700 ;
        RECT 122.460 34.960 122.630 44.050 ;
        RECT 123.245 43.540 123.575 43.710 ;
        RECT 123.030 35.685 123.200 43.325 ;
        RECT 123.620 35.685 123.790 43.325 ;
        RECT 123.245 35.300 123.575 35.470 ;
        RECT 124.190 34.960 124.360 44.050 ;
        RECT 122.460 34.950 124.360 34.960 ;
        RECT 129.460 44.050 131.360 44.220 ;
        RECT 122.290 34.400 124.540 34.950 ;
        RECT 129.460 34.600 129.630 44.050 ;
        RECT 130.245 43.540 130.575 43.710 ;
        RECT 130.030 35.285 130.200 43.325 ;
        RECT 130.620 35.285 130.790 43.325 ;
        RECT 130.245 34.900 130.575 35.070 ;
        RECT 131.190 34.600 131.360 44.050 ;
        RECT 129.240 34.100 131.590 34.600 ;
        RECT 133.060 27.250 133.230 44.600 ;
        RECT 133.845 44.090 134.175 44.260 ;
        RECT 133.630 27.835 133.800 43.875 ;
        RECT 134.220 27.835 134.390 43.875 ;
        RECT 133.845 27.450 134.175 27.620 ;
        RECT 134.790 27.250 134.960 44.600 ;
        RECT 132.840 26.800 135.190 27.250 ;
      LAYER met1 ;
        RECT 103.140 95.450 104.140 96.450 ;
        RECT 104.890 95.400 105.890 96.400 ;
        RECT 112.940 95.400 113.940 96.400 ;
        RECT 114.490 95.350 115.490 96.350 ;
        RECT 126.590 95.400 128.240 96.950 ;
        RECT 0.000 91.750 3.000 92.000 ;
        RECT 98.340 91.750 135.440 94.850 ;
        RECT 0.000 91.150 135.440 91.750 ;
        RECT 0.000 80.600 112.740 91.150 ;
        RECT 122.440 83.850 131.690 91.150 ;
        RECT 133.040 90.300 135.390 91.150 ;
        RECT 133.990 89.900 134.390 90.150 ;
        RECT 134.590 89.695 134.940 90.300 ;
        RECT 122.440 82.600 124.690 83.850 ;
        RECT 129.290 82.950 131.640 83.850 ;
        RECT 123.390 82.050 123.740 82.350 ;
        RECT 123.940 81.845 124.140 82.600 ;
        RECT 130.290 82.400 130.640 82.750 ;
        RECT 130.840 82.245 131.140 82.950 ;
        RECT 0.000 80.250 3.000 80.600 ;
        RECT 100.040 79.500 112.740 80.600 ;
        RECT 100.090 79.000 102.740 79.500 ;
        RECT 101.240 78.450 101.640 78.750 ;
        RECT 101.840 78.265 102.190 79.000 ;
        RECT 100.960 77.950 101.190 78.265 ;
        RECT 100.690 77.265 101.190 77.950 ;
        RECT 101.650 77.600 102.190 78.265 ;
        RECT 101.650 77.265 101.880 77.600 ;
        RECT 103.040 77.550 104.140 78.600 ;
        RECT 110.190 78.500 112.590 79.500 ;
        RECT 111.240 77.950 111.590 78.250 ;
        RECT 111.265 77.900 111.555 77.950 ;
        RECT 111.790 77.695 112.040 78.500 ;
        RECT 103.040 77.500 104.040 77.550 ;
        RECT 100.690 76.250 101.040 77.265 ;
        RECT 101.240 77.050 101.600 77.060 ;
        RECT 103.040 77.050 103.490 77.500 ;
        RECT 111.000 77.400 111.230 77.695 ;
        RECT 101.240 76.750 103.490 77.050 ;
        RECT 110.740 76.695 111.230 77.400 ;
        RECT 111.590 77.150 112.040 77.695 ;
        RECT 111.590 76.695 111.820 77.150 ;
        RECT 112.990 76.850 113.990 77.050 ;
        RECT 100.690 75.900 102.190 76.250 ;
        RECT 101.240 74.850 101.640 75.150 ;
        RECT 101.840 74.685 102.190 75.900 ;
        RECT 110.740 75.700 111.040 76.695 ;
        RECT 112.690 76.550 113.990 76.850 ;
        RECT 111.240 76.200 113.990 76.550 ;
        RECT 112.690 75.850 113.990 76.200 ;
        RECT 112.990 75.750 113.990 75.850 ;
        RECT 110.740 75.400 112.090 75.700 ;
        RECT 100.980 74.200 101.210 74.685 ;
        RECT 100.790 73.685 101.210 74.200 ;
        RECT 101.670 74.200 102.190 74.685 ;
        RECT 111.240 74.650 111.590 74.950 ;
        RECT 111.790 74.445 112.090 75.400 ;
        RECT 123.150 74.900 123.380 81.845 ;
        RECT 101.670 73.685 101.900 74.200 ;
        RECT 111.000 73.950 111.230 74.445 ;
        RECT 98.740 72.500 99.840 72.700 ;
        RECT 100.790 72.500 101.040 73.685 ;
        RECT 98.740 71.500 101.040 72.500 ;
        RECT 98.740 71.150 99.840 71.500 ;
        RECT 100.790 70.460 101.040 71.500 ;
        RECT 101.240 72.500 101.690 73.500 ;
        RECT 110.840 73.445 111.230 73.950 ;
        RECT 111.590 73.900 112.090 74.445 ;
        RECT 122.940 74.245 123.380 74.900 ;
        RECT 123.740 81.350 124.140 81.845 ;
        RECT 123.740 74.245 123.970 81.350 ;
        RECT 130.050 75.200 130.280 82.245 ;
        RECT 129.790 74.245 130.280 75.200 ;
        RECT 130.640 81.550 131.140 82.245 ;
        RECT 130.640 74.245 130.870 81.550 ;
        RECT 111.590 73.445 111.820 73.900 ;
        RECT 108.440 72.550 109.540 72.850 ;
        RECT 101.240 72.300 103.840 72.500 ;
        RECT 101.240 72.150 107.690 72.300 ;
        RECT 108.440 72.200 110.290 72.550 ;
        RECT 110.840 72.200 111.040 73.445 ;
        RECT 101.240 71.600 107.740 72.150 ;
        RECT 101.240 71.500 103.840 71.600 ;
        RECT 101.240 70.600 101.690 71.500 ;
        RECT 100.790 70.050 101.240 70.460 ;
        RECT 101.010 69.960 101.240 70.050 ;
        RECT 101.700 70.200 101.930 70.460 ;
        RECT 101.700 69.960 102.140 70.200 ;
        RECT 101.240 69.550 101.690 69.800 ;
        RECT 101.890 68.950 102.140 69.960 ;
        RECT 100.790 68.750 102.140 68.950 ;
        RECT 100.790 67.700 101.040 68.750 ;
        RECT 106.540 68.350 107.740 71.600 ;
        RECT 108.440 71.800 111.040 72.200 ;
        RECT 108.440 71.550 110.290 71.800 ;
        RECT 108.440 71.300 109.540 71.550 ;
        RECT 110.840 70.700 111.040 71.800 ;
        RECT 111.240 72.200 111.590 73.300 ;
        RECT 119.990 72.550 121.840 73.300 ;
        RECT 122.940 72.550 123.190 74.245 ;
        RECT 112.590 72.200 117.140 72.550 ;
        RECT 111.240 71.800 117.140 72.200 ;
        RECT 111.240 70.850 111.590 71.800 ;
        RECT 112.590 71.750 117.140 71.800 ;
        RECT 112.590 71.550 113.590 71.750 ;
        RECT 110.840 70.200 111.230 70.700 ;
        RECT 111.590 70.550 111.820 70.700 ;
        RECT 111.590 70.200 112.040 70.550 ;
        RECT 111.240 69.800 111.590 70.050 ;
        RECT 111.790 69.400 112.040 70.200 ;
        RECT 116.240 69.950 117.140 71.750 ;
        RECT 119.990 71.550 123.190 72.550 ;
        RECT 119.990 70.950 121.840 71.550 ;
        RECT 110.790 69.150 112.040 69.400 ;
        RECT 112.590 69.450 113.590 69.500 ;
        RECT 114.390 69.450 115.490 69.950 ;
        RECT 101.240 67.850 105.890 68.100 ;
        RECT 100.790 67.450 101.250 67.700 ;
        RECT 101.020 67.200 101.250 67.450 ;
        RECT 101.710 67.500 101.940 67.700 ;
        RECT 101.710 67.200 102.140 67.500 ;
        RECT 101.240 66.800 101.690 67.050 ;
        RECT 101.840 66.500 102.140 67.200 ;
        RECT 102.840 67.150 105.890 67.850 ;
        RECT 110.790 67.650 111.040 69.150 ;
        RECT 112.590 68.850 115.490 69.450 ;
        RECT 111.240 68.650 115.490 68.850 ;
        RECT 111.240 68.500 113.590 68.650 ;
        RECT 111.240 68.040 111.590 68.500 ;
        RECT 114.390 68.350 115.490 68.650 ;
        RECT 116.040 68.300 117.290 69.950 ;
        RECT 122.940 69.500 123.190 71.550 ;
        RECT 123.390 72.550 123.740 74.050 ;
        RECT 125.990 72.550 127.740 72.750 ;
        RECT 129.790 72.550 130.090 74.245 ;
        RECT 130.315 74.000 130.605 74.040 ;
        RECT 133.800 74.000 134.030 89.695 ;
        RECT 130.290 72.550 130.640 74.000 ;
        RECT 133.640 73.695 134.030 74.000 ;
        RECT 134.390 89.250 134.940 89.695 ;
        RECT 134.390 73.695 134.620 89.250 ;
        RECT 123.390 72.350 133.040 72.550 ;
        RECT 133.640 72.350 133.840 73.695 ;
        RECT 134.065 73.400 134.355 73.490 ;
        RECT 123.390 71.900 133.840 72.350 ;
        RECT 123.390 71.550 133.040 71.900 ;
        RECT 123.390 69.650 123.740 71.550 ;
        RECT 125.990 70.450 127.740 71.550 ;
        RECT 122.940 68.950 123.380 69.500 ;
        RECT 111.215 67.810 111.590 68.040 ;
        RECT 111.240 67.800 111.590 67.810 ;
        RECT 110.790 67.350 111.180 67.650 ;
        RECT 110.950 67.150 111.180 67.350 ;
        RECT 111.540 67.500 111.770 67.650 ;
        RECT 111.540 67.150 112.040 67.500 ;
        RECT 102.840 66.900 103.840 67.150 ;
        RECT 111.240 66.990 111.590 67.000 ;
        RECT 111.215 66.760 111.590 66.990 ;
        RECT 111.240 66.750 111.590 66.760 ;
        RECT 100.290 66.100 102.640 66.500 ;
        RECT 111.740 66.450 112.040 67.150 ;
        RECT 110.240 66.100 112.640 66.450 ;
        RECT 100.290 65.050 112.790 66.100 ;
        RECT 123.150 65.700 123.380 68.950 ;
        RECT 123.740 66.150 123.970 69.500 ;
        RECT 129.790 69.450 130.090 71.550 ;
        RECT 130.290 69.600 130.640 71.550 ;
        RECT 133.640 70.650 133.840 71.900 ;
        RECT 134.040 72.350 134.390 73.400 ;
        RECT 136.250 72.700 137.950 73.350 ;
        RECT 135.990 72.550 137.950 72.700 ;
        RECT 135.140 72.350 137.950 72.550 ;
        RECT 134.040 71.900 137.950 72.350 ;
        RECT 134.040 71.200 134.390 71.900 ;
        RECT 135.140 71.550 137.950 71.900 ;
        RECT 135.990 71.400 137.950 71.550 ;
        RECT 135.990 71.300 137.640 71.400 ;
        RECT 134.040 70.800 134.440 71.200 ;
        RECT 133.640 70.200 134.030 70.650 ;
        RECT 129.790 68.700 130.280 69.450 ;
        RECT 123.740 65.700 124.240 66.150 ;
        RECT 123.390 65.250 123.740 65.550 ;
        RECT 3.700 61.500 6.700 61.700 ;
        RECT 100.390 61.550 112.790 65.050 ;
        RECT 123.940 65.000 124.240 65.700 ;
        RECT 130.050 65.450 130.280 68.700 ;
        RECT 130.640 66.250 130.870 69.450 ;
        RECT 130.640 65.450 131.140 66.250 ;
        RECT 122.390 64.200 124.690 65.000 ;
        RECT 130.290 64.950 130.640 65.300 ;
        RECT 130.840 64.750 131.140 65.450 ;
        RECT 129.290 64.200 131.590 64.750 ;
        RECT 122.240 61.550 131.690 64.200 ;
        RECT 133.800 62.650 134.030 70.200 ;
        RECT 134.390 63.080 134.620 70.650 ;
        RECT 134.390 62.650 134.830 63.080 ;
        RECT 134.065 62.460 134.355 62.490 ;
        RECT 134.050 62.120 134.390 62.460 ;
        RECT 134.620 61.900 134.830 62.650 ;
        RECT 133.040 61.550 135.340 61.900 ;
        RECT 98.390 61.500 135.340 61.550 ;
        RECT 3.700 56.000 135.340 61.500 ;
        RECT 3.700 55.900 99.350 56.000 ;
        RECT 3.700 55.700 6.700 55.900 ;
        RECT 100.390 53.300 112.790 56.000 ;
        RECT 100.290 52.750 112.790 53.300 ;
        RECT 122.240 53.550 131.690 56.000 ;
        RECT 132.840 55.650 135.140 56.000 ;
        RECT 133.850 55.090 134.190 55.430 ;
        RECT 133.865 55.060 134.155 55.090 ;
        RECT 134.420 54.900 134.630 55.650 ;
        RECT 100.290 51.850 102.640 52.750 ;
        RECT 101.240 51.300 101.690 51.550 ;
        RECT 101.840 51.150 102.140 51.850 ;
        RECT 110.140 51.750 112.540 52.750 ;
        RECT 122.240 52.550 124.540 53.550 ;
        RECT 129.240 52.800 131.540 53.550 ;
        RECT 123.240 52.000 123.590 52.300 ;
        RECT 123.790 51.850 124.090 52.550 ;
        RECT 130.240 52.250 130.590 52.600 ;
        RECT 130.790 52.100 131.090 52.800 ;
        RECT 101.020 50.900 101.250 51.150 ;
        RECT 100.790 50.650 101.250 50.900 ;
        RECT 101.710 50.850 102.140 51.150 ;
        RECT 102.840 51.100 103.840 51.450 ;
        RECT 111.140 51.440 111.490 51.450 ;
        RECT 104.840 51.100 106.090 51.400 ;
        RECT 111.115 51.210 111.490 51.440 ;
        RECT 111.140 51.200 111.490 51.210 ;
        RECT 101.710 50.650 101.940 50.850 ;
        RECT 100.790 49.600 101.040 50.650 ;
        RECT 102.840 50.500 106.090 51.100 ;
        RECT 111.640 51.050 111.940 51.750 ;
        RECT 110.850 50.850 111.080 51.050 ;
        RECT 101.240 50.300 106.090 50.500 ;
        RECT 110.690 50.550 111.080 50.850 ;
        RECT 111.440 50.700 111.940 51.050 ;
        RECT 111.440 50.550 111.670 50.700 ;
        RECT 101.240 50.250 103.540 50.300 ;
        RECT 104.990 50.200 106.040 50.300 ;
        RECT 100.790 49.400 102.140 49.600 ;
        RECT 101.240 48.550 101.690 48.800 ;
        RECT 101.890 48.390 102.140 49.400 ;
        RECT 101.010 48.300 101.240 48.390 ;
        RECT 100.790 47.890 101.240 48.300 ;
        RECT 101.700 48.150 102.140 48.390 ;
        RECT 106.740 48.350 107.740 49.500 ;
        RECT 110.690 49.050 110.940 50.550 ;
        RECT 111.140 50.390 111.490 50.400 ;
        RECT 111.115 50.160 111.490 50.390 ;
        RECT 111.140 49.700 111.490 50.160 ;
        RECT 113.340 49.700 114.440 49.750 ;
        RECT 111.140 49.350 114.440 49.700 ;
        RECT 110.690 48.800 111.940 49.050 ;
        RECT 101.700 47.890 101.930 48.150 ;
        RECT 98.890 46.850 99.840 47.150 ;
        RECT 100.790 46.850 101.040 47.890 ;
        RECT 98.890 45.850 101.040 46.850 ;
        RECT 98.890 45.700 99.840 45.850 ;
        RECT 100.790 44.665 101.040 45.850 ;
        RECT 101.240 46.850 101.690 47.750 ;
        RECT 106.890 46.850 107.590 48.350 ;
        RECT 111.140 48.150 111.490 48.400 ;
        RECT 111.690 48.000 111.940 48.800 ;
        RECT 112.490 48.700 114.440 49.350 ;
        RECT 115.540 48.250 116.840 49.550 ;
        RECT 123.000 48.600 123.230 51.850 ;
        RECT 110.740 47.500 111.130 48.000 ;
        RECT 111.490 47.650 111.940 48.000 ;
        RECT 111.490 47.500 111.720 47.650 ;
        RECT 101.240 46.150 107.590 46.850 ;
        RECT 101.240 45.850 103.840 46.150 ;
        RECT 106.890 46.100 107.590 46.150 ;
        RECT 108.290 46.650 109.240 47.050 ;
        RECT 108.290 46.400 110.190 46.650 ;
        RECT 110.740 46.400 110.940 47.500 ;
        RECT 108.290 46.000 110.940 46.400 ;
        RECT 101.240 44.850 101.690 45.850 ;
        RECT 108.290 45.650 110.190 46.000 ;
        RECT 108.290 45.600 109.240 45.650 ;
        RECT 110.740 44.755 110.940 46.000 ;
        RECT 111.140 46.400 111.490 47.350 ;
        RECT 115.640 46.750 116.590 48.250 ;
        RECT 122.790 48.050 123.230 48.600 ;
        RECT 123.590 51.400 124.090 51.850 ;
        RECT 123.590 48.050 123.820 51.400 ;
        RECT 130.000 48.850 130.230 52.100 ;
        RECT 129.740 48.100 130.230 48.850 ;
        RECT 130.590 51.300 131.090 52.100 ;
        RECT 130.590 48.100 130.820 51.300 ;
        RECT 113.140 46.650 116.590 46.750 ;
        RECT 112.490 46.400 116.590 46.650 ;
        RECT 111.140 46.000 116.590 46.400 ;
        RECT 111.140 44.900 111.490 46.000 ;
        RECT 112.490 45.650 116.590 46.000 ;
        RECT 119.390 46.000 121.140 47.100 ;
        RECT 122.790 46.000 123.040 48.050 ;
        RECT 119.390 45.000 123.040 46.000 ;
        RECT 119.390 44.800 121.140 45.000 ;
        RECT 100.790 44.150 101.210 44.665 ;
        RECT 100.980 43.665 101.210 44.150 ;
        RECT 101.670 44.150 101.900 44.665 ;
        RECT 110.740 44.250 111.130 44.755 ;
        RECT 101.670 43.665 102.190 44.150 ;
        RECT 110.900 43.755 111.130 44.250 ;
        RECT 111.490 44.300 111.720 44.755 ;
        RECT 111.490 43.755 111.990 44.300 ;
        RECT 101.240 43.200 101.640 43.500 ;
        RECT 101.840 42.450 102.190 43.665 ;
        RECT 111.140 43.250 111.490 43.550 ;
        RECT 111.690 42.800 111.990 43.755 ;
        RECT 100.690 42.100 102.190 42.450 ;
        RECT 110.640 42.500 111.990 42.800 ;
        RECT 122.790 43.305 123.040 45.000 ;
        RECT 123.240 46.000 123.590 47.900 ;
        RECT 126.040 46.000 127.890 47.350 ;
        RECT 129.740 46.000 130.040 48.100 ;
        RECT 130.240 46.000 130.590 47.950 ;
        RECT 133.600 47.350 133.830 54.900 ;
        RECT 133.440 46.900 133.830 47.350 ;
        RECT 134.190 54.470 134.630 54.900 ;
        RECT 134.190 46.900 134.420 54.470 ;
        RECT 123.240 45.650 132.840 46.000 ;
        RECT 133.440 45.650 133.640 46.900 ;
        RECT 123.240 45.200 133.640 45.650 ;
        RECT 123.240 45.000 132.840 45.200 ;
        RECT 123.240 43.500 123.590 45.000 ;
        RECT 129.740 43.305 130.040 45.000 ;
        RECT 130.240 43.550 130.590 45.000 ;
        RECT 133.440 43.855 133.640 45.200 ;
        RECT 133.840 46.350 134.240 46.750 ;
        RECT 133.840 45.650 134.190 46.350 ;
        RECT 135.900 46.250 139.550 46.700 ;
        RECT 135.640 46.000 139.550 46.250 ;
        RECT 134.940 45.650 139.550 46.000 ;
        RECT 133.840 45.200 139.550 45.650 ;
        RECT 133.840 44.150 134.190 45.200 ;
        RECT 134.940 45.000 139.550 45.200 ;
        RECT 135.640 44.850 139.550 45.000 ;
        RECT 135.900 44.700 139.550 44.850 ;
        RECT 133.865 44.060 134.155 44.150 ;
        RECT 133.440 43.550 133.830 43.855 ;
        RECT 130.265 43.510 130.555 43.550 ;
        RECT 122.790 42.650 123.230 43.305 ;
        RECT 100.690 41.085 101.040 42.100 ;
        RECT 101.240 41.300 103.490 41.600 ;
        RECT 101.240 41.290 101.600 41.300 ;
        RECT 103.040 41.200 103.490 41.300 ;
        RECT 110.640 41.505 110.940 42.500 ;
        RECT 113.090 42.350 114.290 42.400 ;
        RECT 112.590 42.000 114.290 42.350 ;
        RECT 111.140 41.650 114.290 42.000 ;
        RECT 100.690 40.400 101.190 41.085 ;
        RECT 100.960 40.085 101.190 40.400 ;
        RECT 101.650 40.750 101.880 41.085 ;
        RECT 101.650 40.085 102.190 40.750 ;
        RECT 101.240 39.600 101.640 39.900 ;
        RECT 101.840 39.350 102.190 40.085 ;
        RECT 103.040 39.850 104.290 41.200 ;
        RECT 110.640 40.800 111.130 41.505 ;
        RECT 110.900 40.505 111.130 40.800 ;
        RECT 111.490 41.050 111.720 41.505 ;
        RECT 112.590 41.350 114.290 41.650 ;
        RECT 111.490 40.505 111.940 41.050 ;
        RECT 113.090 41.000 114.290 41.350 ;
        RECT 111.165 40.250 111.455 40.300 ;
        RECT 111.140 39.950 111.490 40.250 ;
        RECT 111.690 39.700 111.940 40.505 ;
        RECT 100.090 38.800 102.740 39.350 ;
        RECT 110.090 38.800 112.490 39.700 ;
        RECT 0.000 35.700 3.000 35.950 ;
        RECT 100.040 35.700 112.490 38.800 ;
        RECT 123.000 35.705 123.230 42.650 ;
        RECT 123.590 36.200 123.820 43.305 ;
        RECT 129.740 42.350 130.230 43.305 ;
        RECT 123.590 35.705 123.990 36.200 ;
        RECT 0.000 26.300 112.490 35.700 ;
        RECT 123.240 35.200 123.590 35.500 ;
        RECT 123.790 34.950 123.990 35.705 ;
        RECT 130.000 35.305 130.230 42.350 ;
        RECT 130.590 36.000 130.820 43.305 ;
        RECT 130.590 35.305 131.090 36.000 ;
        RECT 122.290 34.150 124.540 34.950 ;
        RECT 130.240 34.800 130.590 35.150 ;
        RECT 130.790 34.600 131.090 35.305 ;
        RECT 129.240 34.150 131.590 34.600 ;
        RECT 122.290 33.400 131.740 34.150 ;
        RECT 122.540 26.300 131.740 33.400 ;
        RECT 133.600 27.855 133.830 43.550 ;
        RECT 134.190 28.300 134.420 43.855 ;
        RECT 134.190 27.855 134.740 28.300 ;
        RECT 133.790 27.400 134.190 27.650 ;
        RECT 134.390 27.250 134.740 27.855 ;
        RECT 132.840 26.300 135.190 27.250 ;
        RECT 0.000 24.550 135.440 26.300 ;
        RECT 0.000 24.400 3.000 24.550 ;
        RECT 98.390 22.850 135.440 24.550 ;
        RECT 103.590 21.300 104.590 22.300 ;
        RECT 105.090 21.400 106.090 22.400 ;
        RECT 113.190 21.300 114.190 22.300 ;
        RECT 115.990 21.000 117.340 22.350 ;
        RECT 125.800 19.850 128.500 21.550 ;
        RECT 126.140 19.800 128.390 19.850 ;
      LAYER met2 ;
        RECT 102.800 95.350 104.150 96.600 ;
        RECT 104.750 95.400 105.950 96.600 ;
        RECT 0.000 80.250 3.000 92.000 ;
        RECT 103.090 78.600 104.140 95.350 ;
        RECT 103.040 77.550 104.140 78.600 ;
        RECT 98.740 71.150 99.840 72.700 ;
        RECT 98.890 64.250 99.740 71.150 ;
        RECT 104.840 67.150 105.890 95.400 ;
        RECT 112.750 95.350 113.940 96.540 ;
        RECT 114.450 95.350 115.550 96.550 ;
        RECT 126.200 95.400 128.400 97.050 ;
        RECT 113.240 77.050 113.940 95.350 ;
        RECT 112.990 75.750 113.990 77.050 ;
        RECT 108.440 71.300 109.540 72.850 ;
        RECT 106.590 68.450 107.690 70.050 ;
        RECT 108.540 64.250 109.390 71.300 ;
        RECT 114.490 69.950 115.340 95.350 ;
        RECT 117.790 75.500 119.390 75.550 ;
        RECT 126.590 75.500 128.240 95.400 ;
        RECT 117.740 74.500 128.240 75.500 ;
        RECT 117.740 73.800 127.690 74.500 ;
        RECT 114.390 68.350 115.490 69.950 ;
        RECT 116.040 68.300 117.290 69.950 ;
        RECT 98.890 63.850 116.440 64.250 ;
        RECT 98.940 63.150 116.440 63.850 ;
        RECT 3.700 61.500 6.700 61.700 ;
        RECT 3.700 61.495 9.300 61.500 ;
        RECT 3.700 55.905 92.445 61.495 ;
        RECT 3.700 55.900 9.300 55.905 ;
        RECT 3.700 55.700 6.700 55.900 ;
        RECT 117.790 54.950 119.390 73.800 ;
        RECT 119.990 70.950 121.840 73.300 ;
        RECT 126.190 72.750 127.690 73.800 ;
        RECT 125.990 71.400 127.740 72.750 ;
        RECT 120.190 60.650 121.540 70.950 ;
        RECT 125.990 70.450 127.840 71.400 ;
        RECT 126.240 68.300 127.840 70.450 ;
        RECT 120.190 60.400 127.540 60.650 ;
        RECT 120.190 58.750 127.640 60.400 ;
        RECT 120.190 58.700 121.540 58.750 ;
        RECT 98.390 53.900 119.390 54.950 ;
        RECT 98.390 47.150 99.140 53.900 ;
        RECT 104.840 50.200 106.090 51.350 ;
        RECT 98.390 46.450 99.840 47.150 ;
        RECT 98.890 45.700 99.840 46.450 ;
        RECT 103.040 40.800 104.290 41.200 ;
        RECT 103.040 39.850 104.340 40.800 ;
        RECT 0.000 24.400 3.000 35.950 ;
        RECT 103.640 22.500 104.340 39.850 ;
        RECT 105.140 22.500 105.940 50.200 ;
        RECT 106.740 48.350 107.740 49.500 ;
        RECT 108.290 47.050 109.040 53.900 ;
        RECT 113.340 48.700 114.440 49.750 ;
        RECT 108.290 45.600 109.240 47.050 ;
        RECT 113.540 44.100 114.440 48.700 ;
        RECT 115.540 48.250 116.940 49.500 ;
        RECT 117.790 47.100 119.390 53.900 ;
        RECT 126.290 49.600 127.640 58.750 ;
        RECT 126.190 48.350 127.640 49.600 ;
        RECT 126.290 47.350 127.640 48.350 ;
        RECT 126.040 47.250 127.890 47.350 ;
        RECT 117.790 44.850 121.140 47.100 ;
        RECT 126.040 45.000 128.390 47.250 ;
        RECT 119.390 44.800 121.140 44.850 ;
        RECT 113.540 43.350 117.190 44.100 ;
        RECT 103.150 20.900 104.600 22.500 ;
        RECT 105.050 20.900 106.500 22.500 ;
        RECT 113.090 22.330 114.290 42.400 ;
        RECT 116.290 22.400 117.190 43.350 ;
        RECT 112.500 20.500 114.290 22.330 ;
        RECT 115.800 20.350 117.450 22.400 ;
        RECT 126.140 21.650 128.390 45.000 ;
        RECT 130.690 26.200 133.390 94.350 ;
        RECT 151.350 73.200 153.000 73.350 ;
        RECT 136.400 71.250 153.000 73.200 ;
        RECT 151.350 71.050 153.000 71.250 ;
        RECT 135.900 44.700 139.550 46.700 ;
        RECT 130.490 22.950 133.390 26.200 ;
        RECT 125.650 19.500 128.600 21.650 ;
      LAYER met3 ;
        RECT 100.550 215.300 119.575 216.450 ;
        RECT 104.750 213.155 122.420 214.300 ;
        RECT 104.750 213.150 106.000 213.155 ;
        RECT 116.050 209.200 125.125 210.350 ;
        RECT 114.200 207.250 127.875 208.400 ;
        RECT 96.825 204.200 130.550 205.350 ;
        RECT 102.825 202.100 133.400 203.250 ;
        RECT 110.525 199.600 136.050 200.750 ;
        RECT 112.775 197.350 138.900 198.500 ;
        RECT 102.800 95.350 104.150 96.600 ;
        RECT 104.750 95.400 105.950 96.600 ;
        RECT 112.750 95.350 113.940 96.540 ;
        RECT 114.450 95.350 115.550 96.550 ;
        RECT 126.200 95.400 128.400 97.050 ;
        RECT 0.000 80.250 3.000 92.000 ;
        RECT 151.350 71.050 153.000 73.350 ;
        RECT 106.740 68.400 127.890 69.750 ;
        RECT 115.040 62.950 121.590 64.550 ;
        RECT 3.700 55.700 6.700 61.700 ;
        RECT 106.740 49.350 107.740 49.500 ;
        RECT 126.190 49.350 127.590 49.600 ;
        RECT 106.740 48.400 127.590 49.350 ;
        RECT 106.740 48.350 107.740 48.400 ;
        RECT 126.190 48.350 127.590 48.400 ;
        RECT 135.900 44.700 139.550 46.700 ;
        RECT 0.000 24.400 3.000 35.950 ;
        RECT 103.150 20.900 104.600 22.500 ;
        RECT 105.050 20.900 106.500 22.500 ;
        RECT 112.500 20.500 114.290 22.330 ;
        RECT 115.800 20.350 117.450 22.400 ;
        RECT 125.650 19.500 128.600 21.650 ;
      LAYER met4 ;
        RECT 121.600 224.760 121.750 224.795 ;
        RECT 122.050 224.760 122.250 224.795 ;
        RECT 100.550 215.300 101.800 216.450 ;
        RECT 0.000 80.250 1.000 92.000 ;
        RECT 3.700 55.700 4.000 61.700 ;
        RECT 6.000 55.700 6.700 61.700 ;
        RECT 0.000 24.400 1.000 35.950 ;
        RECT 97.215 25.435 98.185 205.885 ;
        RECT 100.655 93.960 101.645 215.300 ;
        RECT 118.785 215.225 119.435 224.760 ;
        RECT 104.750 213.150 106.000 214.300 ;
        RECT 102.960 98.700 103.990 203.500 ;
        RECT 102.950 96.600 104.000 98.700 ;
        RECT 104.850 96.600 105.900 213.150 ;
        RECT 121.600 212.775 122.250 224.760 ;
        RECT 124.345 224.760 124.510 224.855 ;
        RECT 124.810 224.760 124.995 224.855 ;
        RECT 116.050 209.200 117.300 210.350 ;
        RECT 114.200 207.250 115.450 208.400 ;
        RECT 102.800 95.350 104.150 96.600 ;
        RECT 104.750 95.400 105.950 96.600 ;
        RECT 100.640 92.935 106.240 93.960 ;
        RECT 105.215 25.650 106.240 92.935 ;
        RECT 110.755 91.890 111.945 201.050 ;
        RECT 112.915 103.050 113.790 198.650 ;
        RECT 112.900 96.540 113.800 103.050 ;
        RECT 114.550 96.550 115.450 207.250 ;
        RECT 112.750 95.350 113.940 96.540 ;
        RECT 114.450 95.350 115.550 96.550 ;
        RECT 110.755 90.705 115.090 91.890 ;
        RECT 110.755 90.700 111.945 90.705 ;
        RECT 113.905 29.775 115.090 90.705 ;
        RECT 112.925 28.605 115.090 29.775 ;
        RECT 112.925 26.300 114.080 28.605 ;
        RECT 101.385 25.435 104.415 25.465 ;
        RECT 97.215 24.465 104.415 25.435 ;
        RECT 101.385 24.435 104.415 24.465 ;
        RECT 103.385 22.500 104.415 24.435 ;
        RECT 105.200 22.500 106.250 25.650 ;
        RECT 103.150 20.900 104.600 22.500 ;
        RECT 105.050 20.900 106.500 22.500 ;
        RECT 112.900 22.330 114.100 26.300 ;
        RECT 116.105 25.750 117.300 209.200 ;
        RECT 124.345 208.875 124.995 224.760 ;
        RECT 127.095 224.760 127.270 224.855 ;
        RECT 127.570 224.760 127.745 224.855 ;
        RECT 127.095 206.675 127.745 224.760 ;
        RECT 129.840 224.760 130.030 224.790 ;
        RECT 130.330 224.760 130.490 224.790 ;
        RECT 129.840 205.350 130.490 224.760 ;
        RECT 132.635 224.760 132.790 224.800 ;
        RECT 133.090 224.760 133.285 224.800 ;
        RECT 129.250 204.200 130.550 205.350 ;
        RECT 132.635 203.250 133.285 224.760 ;
        RECT 135.345 224.760 135.550 224.815 ;
        RECT 135.850 224.760 135.995 224.815 ;
        RECT 132.250 202.100 133.400 203.250 ;
        RECT 135.345 200.750 135.995 224.760 ;
        RECT 138.150 224.760 138.310 224.815 ;
        RECT 138.610 224.760 138.800 224.815 ;
        RECT 134.900 199.600 136.050 200.750 ;
        RECT 138.150 198.500 138.800 224.760 ;
        RECT 137.750 197.350 138.900 198.500 ;
        RECT 119.050 97.150 120.350 97.250 ;
        RECT 118.950 97.050 127.900 97.150 ;
        RECT 118.950 95.850 128.400 97.050 ;
        RECT 116.100 22.400 117.300 25.750 ;
        RECT 112.500 20.500 114.290 22.330 ;
        RECT 115.800 20.350 117.450 22.400 ;
        RECT 119.050 16.150 120.350 95.850 ;
        RECT 126.200 95.400 128.400 95.850 ;
        RECT 151.350 71.050 153.000 73.350 ;
        RECT 135.900 46.650 139.550 46.700 ;
        RECT 135.900 44.700 139.650 46.650 ;
        RECT 125.650 19.500 128.600 21.650 ;
        RECT 93.600 14.750 120.350 16.150 ;
        RECT 93.800 1.000 94.800 14.750 ;
        RECT 126.000 12.850 128.300 19.500 ;
        RECT 113.000 11.250 128.300 12.850 ;
        RECT 93.800 0.750 93.850 1.000 ;
        RECT 94.750 0.750 94.800 1.000 ;
        RECT 113.100 1.000 114.100 11.250 ;
        RECT 138.350 10.450 139.650 44.700 ;
        RECT 113.100 0.600 113.170 1.000 ;
        RECT 114.070 0.600 114.100 1.000 ;
        RECT 132.450 8.950 139.650 10.450 ;
        RECT 132.450 1.000 133.400 8.950 ;
        RECT 132.450 0.600 132.490 1.000 ;
        RECT 133.390 0.600 133.400 1.000 ;
        RECT 151.800 1.000 152.800 71.050 ;
        RECT 151.800 0.400 151.810 1.000 ;
        RECT 152.710 0.400 152.800 1.000 ;
  END
END tt_um_sky25a_nurirfansyah_nauta
END LIBRARY

