magic
tech sky130A
magscale 1 2
timestamp 1762798763
<< metal1 >>
rect 200 18350 600 18400
rect 200 16120 250 18350
rect 540 16120 20550 18350
rect 200 16050 600 16120
rect 27250 14600 27590 14670
rect 27250 14330 27280 14600
rect 27520 14330 27590 14600
rect 27250 14280 27590 14330
rect 740 12310 1340 12340
rect 740 11190 790 12310
rect 1300 12300 1340 12310
rect 1300 12130 19870 12300
rect 1300 11380 1640 12130
rect 2610 12110 19870 12130
rect 2610 12090 17230 12110
rect 2610 11380 8780 12090
rect 1300 11340 8780 11380
rect 9750 11360 17230 12090
rect 18200 11360 19870 12110
rect 9750 11340 19870 11360
rect 1300 11190 19870 11340
rect 740 11180 19870 11190
rect 740 11140 1340 11180
rect 27180 9260 27910 9340
rect 27180 9020 27260 9260
rect 27820 9020 27910 9260
rect 27180 8940 27910 9020
rect 200 7140 600 7190
rect 200 4940 250 7140
rect 540 4940 20100 7140
rect 200 4910 20100 4940
rect 200 4880 600 4910
rect 25160 3970 25700 4310
<< via1 >>
rect 250 16120 540 18350
rect 27280 14330 27520 14600
rect 790 11190 1300 12310
rect 1640 11380 2610 12130
rect 8780 11340 9750 12090
rect 17230 11360 18200 12110
rect 27260 9020 27820 9260
rect 250 4940 540 7140
<< metal2 >>
rect 25240 19350 25680 19410
rect 20560 19300 20830 19320
rect 20560 19090 20580 19300
rect 20810 19090 20830 19300
rect 20560 19070 20830 19090
rect 20950 19300 21190 19320
rect 20950 19100 20970 19300
rect 21170 19100 21190 19300
rect 20950 19080 21190 19100
rect 22550 19270 22788 19308
rect 22550 19100 22590 19270
rect 22760 19100 22788 19270
rect 22550 19070 22788 19100
rect 22890 19290 23110 19310
rect 22890 19090 22910 19290
rect 23090 19090 23110 19290
rect 22890 19070 23110 19090
rect 25240 19130 25290 19350
rect 25630 19130 25680 19350
rect 25240 19080 25680 19130
rect 200 18350 600 18400
rect 200 16120 250 18350
rect 540 16120 600 18350
rect 200 16050 600 16120
rect 30270 14640 30600 14670
rect 27280 14600 30290 14640
rect 27520 14330 30290 14600
rect 27280 14280 30290 14330
rect 30530 14280 30600 14640
rect 27280 14250 30600 14280
rect 30270 14210 30600 14250
rect 740 12310 1340 12340
rect 740 11190 790 12310
rect 1300 12300 1340 12310
rect 1300 12299 1860 12300
rect 1300 12130 18489 12299
rect 1300 11380 1640 12130
rect 2610 12110 18489 12130
rect 2610 12090 17230 12110
rect 2610 11380 8780 12090
rect 1300 11340 8780 11380
rect 9750 11360 17230 12090
rect 18200 11360 18489 12110
rect 9750 11340 18489 11360
rect 1300 11190 18489 11340
rect 740 11181 18489 11190
rect 740 11180 1860 11181
rect 740 11140 1340 11180
rect 27180 9260 27910 9340
rect 27180 9020 27260 9260
rect 27820 9020 27910 9260
rect 27180 8940 27910 9020
rect 200 7140 600 7190
rect 200 4940 250 7140
rect 540 4940 600 7140
rect 200 4880 600 4940
rect 20630 4470 20920 4500
rect 20630 4230 20660 4470
rect 20890 4230 20920 4470
rect 20630 4180 20920 4230
rect 21010 4480 21300 4500
rect 21010 4200 21030 4480
rect 21280 4200 21300 4480
rect 21010 4180 21300 4200
rect 22500 4420 22858 4466
rect 22500 4150 22540 4420
rect 22820 4150 22858 4420
rect 22500 4100 22858 4150
rect 23160 4460 23490 4480
rect 23160 4110 23180 4460
rect 23470 4110 23490 4460
rect 23160 4070 23490 4110
rect 25130 4240 25720 4330
rect 25130 3950 25200 4240
rect 25650 3950 25720 4240
rect 25130 3900 25720 3950
<< via2 >>
rect 20580 19090 20810 19300
rect 20970 19100 21170 19300
rect 22590 19100 22760 19270
rect 22910 19090 23090 19290
rect 25290 19130 25630 19350
rect 250 16120 540 18350
rect 30290 14280 30530 14640
rect 790 11190 1300 12310
rect 27260 9020 27820 9260
rect 250 4940 540 7140
rect 20660 4230 20890 4470
rect 21030 4200 21280 4480
rect 22540 4150 22820 4420
rect 23180 4110 23470 4460
rect 25200 3950 25650 4240
<< metal3 >>
rect 20110 43270 23915 43290
rect 20110 43090 20130 43270
rect 20340 43260 23915 43270
rect 20340 43090 23770 43260
rect 20110 43080 23770 43090
rect 23870 43080 23915 43260
rect 20110 43060 23915 43080
rect 20950 42840 24484 42860
rect 20950 42670 20970 42840
rect 21170 42670 24330 42840
rect 20950 42660 24330 42670
rect 24430 42660 24484 42840
rect 20950 42631 24484 42660
rect 20950 42630 21200 42631
rect 23210 42050 25025 42070
rect 23210 42040 24880 42050
rect 23210 41870 23250 42040
rect 23430 41870 24880 42040
rect 23210 41860 24880 41870
rect 24980 41860 25025 42050
rect 23210 41840 25025 41860
rect 22840 41660 25575 41680
rect 22840 41650 25430 41660
rect 22840 41480 22870 41650
rect 23050 41480 25430 41650
rect 22840 41470 25430 41480
rect 25530 41470 25575 41660
rect 22840 41450 25575 41470
rect 19365 41050 26110 41070
rect 19365 40860 19460 41050
rect 19620 40860 25880 41050
rect 26080 40860 26110 41050
rect 19365 40840 26110 40860
rect 20565 40630 26680 40650
rect 20565 40440 20610 40630
rect 20780 40440 26470 40630
rect 26660 40440 26680 40630
rect 20565 40420 26680 40440
rect 22105 40130 27210 40150
rect 22105 39940 22170 40130
rect 22370 39940 27000 40130
rect 27190 39940 27210 40130
rect 22105 39920 27210 39940
rect 22555 39680 27780 39700
rect 22555 39490 22610 39680
rect 22740 39490 27570 39680
rect 27760 39490 27780 39680
rect 22555 39470 27780 39490
rect 25240 19350 25680 19410
rect 20560 19300 20830 19320
rect 20560 19090 20580 19300
rect 20810 19090 20830 19300
rect 20560 19070 20830 19090
rect 20950 19300 21190 19320
rect 20950 19100 20970 19300
rect 21170 19100 21190 19300
rect 20950 19080 21190 19100
rect 22550 19270 22788 19308
rect 22550 19100 22590 19270
rect 22760 19100 22788 19270
rect 22550 19070 22788 19100
rect 22890 19290 23110 19310
rect 22890 19090 22910 19290
rect 23090 19090 23110 19290
rect 22890 19070 23110 19090
rect 25240 19130 25290 19350
rect 25630 19130 25680 19350
rect 25240 19080 25680 19130
rect 200 18350 600 18400
rect 200 16120 250 18350
rect 540 16120 600 18350
rect 200 16050 600 16120
rect 30270 14640 30600 14670
rect 30270 14280 30290 14640
rect 30530 14280 30600 14640
rect 30270 14210 30600 14280
rect 740 12310 1340 12340
rect 740 11190 790 12310
rect 1300 11190 1340 12310
rect 740 11140 1340 11190
rect 27180 9260 27910 9340
rect 27180 9020 27260 9260
rect 27820 9020 27910 9260
rect 27180 8940 27910 9020
rect 200 7140 600 7190
rect 200 4940 250 7140
rect 540 4940 600 7140
rect 200 4880 600 4940
rect 20630 4470 20920 4500
rect 20630 4230 20660 4470
rect 20890 4230 20920 4470
rect 20630 4180 20920 4230
rect 21010 4480 21300 4500
rect 21010 4200 21030 4480
rect 21280 4200 21300 4480
rect 21010 4180 21300 4200
rect 22500 4420 22858 4466
rect 22500 4150 22540 4420
rect 22820 4150 22858 4420
rect 22500 4100 22858 4150
rect 23160 4460 23490 4480
rect 23160 4110 23180 4460
rect 23470 4110 23490 4460
rect 23160 4070 23490 4110
rect 25130 4240 25720 4330
rect 25130 3950 25200 4240
rect 25650 3950 25720 4240
rect 25130 3900 25720 3950
<< via3 >>
rect 20130 43090 20340 43270
rect 23770 43080 23870 43260
rect 20970 42670 21170 42840
rect 24330 42660 24430 42840
rect 23250 41870 23430 42040
rect 24880 41860 24980 42050
rect 22870 41480 23050 41650
rect 25430 41470 25530 41660
rect 19460 40860 19620 41050
rect 25880 40860 26080 41050
rect 20610 40440 20780 40630
rect 26470 40440 26660 40630
rect 22170 39940 22370 40130
rect 27000 39940 27190 40130
rect 22610 39490 22740 39680
rect 27570 39490 27760 39680
rect 20580 19090 20810 19300
rect 20970 19100 21170 19300
rect 22590 19100 22760 19270
rect 22910 19090 23090 19290
rect 25290 19130 25630 19350
rect 250 16120 540 18350
rect 30290 14280 30530 14640
rect 790 11190 1300 12310
rect 27260 9020 27820 9260
rect 250 4940 540 7140
rect 20660 4230 20890 4470
rect 21030 4200 21280 4480
rect 22540 4150 22820 4420
rect 23180 4110 23470 4460
rect 25200 3950 25650 4240
<< metal4 >>
rect 6134 44960 6194 45152
rect 6686 44960 6746 45152
rect 7238 44960 7298 45152
rect 7790 44960 7850 45152
rect 8342 44960 8402 45152
rect 8894 44960 8954 45152
rect 9446 44960 9506 45152
rect 9998 44960 10058 45152
rect 10550 44960 10610 45152
rect 11102 44960 11162 45152
rect 11654 44960 11714 45152
rect 12206 44960 12266 45152
rect 12758 44960 12818 45152
rect 13310 44960 13370 45152
rect 13862 44960 13922 45152
rect 14414 44960 14474 45152
rect 14966 44960 15026 45152
rect 15518 44960 15578 45152
rect 16070 44960 16130 45152
rect 16622 44960 16682 45152
rect 17174 44960 17234 45152
rect 17726 44960 17786 45152
rect 18278 44960 18338 45152
rect 18830 44960 18890 45152
rect 6080 44830 18900 44960
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44959 24410 45152
rect 24902 44971 24962 45152
rect 25454 44971 25514 45152
rect 200 18350 600 44152
rect 200 16120 250 18350
rect 540 16120 600 18350
rect 200 7140 600 16120
rect 800 43980 1200 44152
rect 7390 43980 7580 44830
rect 800 43700 7580 43980
rect 800 12340 1200 43700
rect 20110 43270 20360 43290
rect 20110 43090 20130 43270
rect 20340 43090 20360 43270
rect 20110 43060 20360 43090
rect 23757 43260 23887 44952
rect 23757 43080 23770 43260
rect 23870 43080 23887 43260
rect 19443 41050 19637 41177
rect 19443 40860 19460 41050
rect 19620 40860 19637 41050
rect 740 12310 1340 12340
rect 740 11190 790 12310
rect 1300 11190 1340 12310
rect 740 11140 1340 11190
rect 200 4940 250 7140
rect 540 4940 600 7140
rect 200 1000 600 4940
rect 800 1000 1200 11140
rect 19443 5087 19637 40860
rect 20131 18792 20329 43060
rect 23757 43045 23887 43080
rect 20950 42840 21200 42860
rect 20950 42670 20970 42840
rect 21170 42670 21200 42840
rect 20950 42630 21200 42670
rect 24320 42840 24450 44959
rect 24320 42660 24330 42840
rect 24430 42660 24450 42840
rect 20592 40630 20798 40700
rect 20592 40440 20610 40630
rect 20780 40440 20798 40630
rect 20592 19740 20798 40440
rect 20590 19320 20800 19740
rect 20970 19320 21180 42630
rect 24320 42555 24450 42660
rect 23210 42040 23460 42070
rect 23210 41870 23250 42040
rect 23430 41870 23460 42040
rect 23210 41840 23460 41870
rect 22840 41650 23090 41680
rect 22840 41480 22870 41650
rect 23050 41480 23090 41650
rect 22840 41450 23090 41480
rect 22151 40130 22389 40210
rect 22151 39940 22170 40130
rect 22370 39940 22389 40130
rect 20560 19300 20830 19320
rect 20560 19090 20580 19300
rect 20810 19090 20830 19300
rect 20560 19070 20830 19090
rect 20950 19300 21190 19320
rect 20950 19100 20970 19300
rect 21170 19100 21190 19300
rect 20950 19080 21190 19100
rect 20128 18587 21248 18792
rect 21043 5130 21248 18587
rect 22151 18378 22389 39940
rect 22583 39680 22758 39730
rect 22583 39490 22610 39680
rect 22740 39490 22758 39680
rect 22583 20610 22758 39490
rect 22580 19308 22760 20610
rect 22910 19310 23090 41450
rect 22550 19270 22788 19308
rect 22550 19100 22590 19270
rect 22760 19100 22788 19270
rect 22550 19070 22788 19100
rect 22890 19290 23110 19310
rect 22890 19090 22910 19290
rect 23090 19090 23110 19290
rect 22890 19070 23110 19090
rect 22151 18141 23018 18378
rect 22151 18140 22389 18141
rect 22781 5955 23018 18141
rect 22585 5721 23018 5955
rect 22585 5260 22816 5721
rect 20277 5087 20883 5093
rect 19443 4893 20883 5087
rect 20277 4887 20883 4893
rect 20677 4500 20883 4887
rect 21040 4500 21250 5130
rect 20630 4470 20920 4500
rect 20630 4230 20660 4470
rect 20890 4230 20920 4470
rect 20630 4180 20920 4230
rect 21010 4480 21300 4500
rect 21010 4200 21030 4480
rect 21280 4200 21300 4480
rect 22580 4466 22820 5260
rect 23221 5150 23460 41840
rect 24869 42050 24999 44971
rect 24869 41860 24880 42050
rect 24980 41860 24999 42050
rect 24869 41775 24999 41860
rect 25419 41660 25549 44971
rect 26006 44958 26066 45152
rect 26558 44960 26618 45152
rect 27110 44963 27170 45152
rect 27662 44963 27722 45152
rect 25419 41470 25430 41660
rect 25530 41470 25549 41660
rect 25419 41335 25549 41470
rect 25968 41070 26098 44958
rect 25850 41050 26110 41070
rect 25850 40860 25880 41050
rect 26080 40860 26110 41050
rect 25850 40840 26110 40860
rect 26527 40650 26657 44960
rect 26450 40630 26680 40650
rect 26450 40440 26470 40630
rect 26660 40440 26680 40630
rect 26450 40420 26680 40440
rect 27069 40150 27199 44963
rect 26980 40130 27210 40150
rect 26980 39940 27000 40130
rect 27190 39940 27210 40130
rect 26980 39920 27210 39940
rect 27630 39700 27760 44963
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27550 39680 27780 39700
rect 27550 39490 27570 39680
rect 27760 39490 27780 39680
rect 27550 39470 27780 39490
rect 23810 19430 24070 19450
rect 23790 19410 25580 19430
rect 23790 19350 25680 19410
rect 23790 19170 25290 19350
rect 23220 4480 23460 5150
rect 21010 4180 21300 4200
rect 22500 4420 22858 4466
rect 22500 4150 22540 4420
rect 22820 4150 22858 4420
rect 22500 4100 22858 4150
rect 23160 4460 23490 4480
rect 23160 4110 23180 4460
rect 23470 4110 23490 4460
rect 23160 4070 23490 4110
rect 23810 3230 24070 19170
rect 25240 19130 25290 19170
rect 25630 19130 25680 19350
rect 25240 19080 25680 19130
rect 30270 14640 30600 14670
rect 30270 14280 30290 14640
rect 30530 14280 30600 14640
rect 30270 14210 30600 14280
rect 27180 9330 27910 9340
rect 27180 9260 27930 9330
rect 27180 9020 27260 9260
rect 27820 9020 27930 9260
rect 27180 8940 27930 9020
rect 25130 4240 25720 4330
rect 25130 3950 25200 4240
rect 25650 3950 25720 4240
rect 25130 3900 25720 3950
rect 18720 2950 24070 3230
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18760 150 18960 2950
rect 25200 2570 25660 3900
rect 22600 2250 25660 2570
rect 18770 0 18950 150
rect 22620 120 22820 2250
rect 27670 2090 27930 8940
rect 26490 1790 27930 2090
rect 26490 120 26680 1790
rect 22634 0 22814 120
rect 26498 0 26678 120
rect 30360 80 30560 14210
rect 30362 0 30542 80
use nauta_ota_dtrim2b  nauta_ota_dtrim2b_0
timestamp 1757964080
transform -1 0 36908 0 1 11000
box 9380 -7040 17240 8390
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
