magic
tech sky130A
magscale 1 2
timestamp 1757958533
<< locali >>
rect 1120 1500 1590 1520
rect 1120 1440 1150 1500
rect 1560 1440 1590 1500
rect 1120 1420 1590 1440
rect 1130 -2240 1590 -2220
rect 1130 -2320 1160 -2240
rect 1560 -2320 1590 -2240
rect 1130 -2340 1590 -2320
<< viali >>
rect 1150 1440 1560 1500
rect 1160 -2320 1560 -2240
<< metal1 >>
rect 1120 1500 1590 1770
rect 1120 1440 1150 1500
rect 1560 1440 1590 1500
rect 1120 1420 1590 1440
rect 1220 1140 1280 1420
rect 1320 1310 1390 1380
rect 1320 -660 1390 -370
rect 1100 -860 1390 -660
rect 1320 -1250 1390 -860
rect 1430 -660 1490 -130
rect 1430 -860 1750 -660
rect 1430 -1430 1490 -860
rect 1220 -2220 1280 -1920
rect 1320 -2180 1390 -2110
rect 1130 -2240 1590 -2220
rect 1130 -2320 1160 -2240
rect 1560 -2320 1590 -2240
rect 1130 -2550 1590 -2320
use sky130_fd_pr__nfet_01v8_SALWK2  XM1
timestamp 1757953701
transform 1 0 1356 0 1 -1680
box -226 -610 226 610
use sky130_fd_pr__pfet_01v8_SKDPWJ  XM2
timestamp 1757953701
transform 1 0 1356 0 1 479
box -226 -1019 226 1019
<< labels >>
flabel metal1 1100 -860 1300 -660 0 FreeSans 256 0 0 0 in
port 1 nsew
flabel metal1 1120 1570 1320 1770 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 1140 -2540 1340 -2340 0 FreeSans 256 0 0 0 gnd
port 3 nsew
flabel metal1 1550 -860 1750 -660 0 FreeSans 256 0 0 0 out
port 2 nsew
<< end >>
