magic
tech sky130A
magscale 1 2
timestamp 1757952087
<< error_p >>
rect -29 872 29 878
rect -29 838 -17 872
rect -29 832 29 838
rect -29 -838 29 -832
rect -29 -872 -17 -838
rect -29 -878 29 -872
<< pwell >>
rect -226 -1010 226 1010
<< nmos >>
rect -30 -800 30 800
<< ndiff >>
rect -88 788 -30 800
rect -88 -788 -76 788
rect -42 -788 -30 788
rect -88 -800 -30 -788
rect 30 788 88 800
rect 30 -788 42 788
rect 76 -788 88 788
rect 30 -800 88 -788
<< ndiffc >>
rect -76 -788 -42 788
rect 42 -788 76 788
<< psubdiff >>
rect -190 940 -94 974
rect 94 940 190 974
rect -190 878 -156 940
rect 156 878 190 940
rect -190 -940 -156 -878
rect 156 -940 190 -878
rect -190 -974 -94 -940
rect 94 -974 190 -940
<< psubdiffcont >>
rect -94 940 94 974
rect -190 -878 -156 878
rect 156 -878 190 878
rect -94 -974 94 -940
<< poly >>
rect -33 872 33 888
rect -33 838 -17 872
rect 17 838 33 872
rect -33 822 33 838
rect -30 800 30 822
rect -30 -822 30 -800
rect -33 -838 33 -822
rect -33 -872 -17 -838
rect 17 -872 33 -838
rect -33 -888 33 -872
<< polycont >>
rect -17 838 17 872
rect -17 -872 17 -838
<< locali >>
rect -190 940 -94 974
rect 94 940 190 974
rect -190 878 -156 940
rect 156 878 190 940
rect -33 838 -17 872
rect 17 838 33 872
rect -76 788 -42 804
rect -76 -804 -42 -788
rect 42 788 76 804
rect 42 -804 76 -788
rect -33 -872 -17 -838
rect 17 -872 33 -838
rect -190 -940 -156 -878
rect 156 -940 190 -878
rect -190 -974 -94 -940
rect 94 -974 190 -940
<< viali >>
rect -17 838 17 872
rect -76 -788 -42 788
rect 42 -788 76 788
rect -17 -872 17 -838
<< metal1 >>
rect -29 872 29 878
rect -29 838 -17 872
rect 17 838 29 872
rect -29 832 29 838
rect -82 788 -36 800
rect -82 -788 -76 788
rect -42 -788 -36 788
rect -82 -800 -36 -788
rect 36 788 82 800
rect 36 -788 42 788
rect 76 -788 82 788
rect 36 -800 82 -788
rect -29 -838 29 -832
rect -29 -872 -17 -838
rect 17 -872 29 -838
rect -29 -878 29 -872
<< properties >>
string FIXED_BBOX -173 -957 173 957
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
