magic
tech sky130A
magscale 1 2
timestamp 1757947919
<< error_p >>
rect -255 997 255 1003
rect -255 969 -249 997
rect 249 969 255 997
rect -255 963 255 969
rect -88 -847 -30 -841
rect 30 -847 88 -841
rect -88 -881 -76 -847
rect 30 -881 42 -847
rect -88 -887 -30 -881
rect 30 -887 88 -881
<< nwell >>
rect -285 -1019 285 1019
<< pmos >>
rect -89 -800 -29 800
rect 29 -800 89 800
<< pdiff >>
rect -147 788 -89 800
rect -147 -788 -135 788
rect -101 -788 -89 788
rect -147 -800 -89 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 89 788 147 800
rect 89 -788 101 788
rect 135 -788 147 788
rect 89 -800 147 -788
<< pdiffc >>
rect -135 -788 -101 788
rect -17 -788 17 788
rect 101 -788 135 788
<< nsubdiff >>
rect -249 949 -153 983
rect 153 949 249 983
rect -249 887 -215 949
rect 215 887 249 949
rect -249 -949 -215 -887
rect 215 -949 249 -887
rect -249 -983 -153 -949
rect 153 -983 249 -949
<< nsubdiffcont >>
rect -153 949 153 983
rect -249 -887 -215 887
rect 215 -887 249 887
rect -153 -983 153 -949
<< poly >>
rect -92 881 -26 897
rect -92 847 -76 881
rect -42 847 -26 881
rect -92 831 -26 847
rect 26 881 92 897
rect 26 847 42 881
rect 76 847 92 881
rect 26 831 92 847
rect -89 800 -29 831
rect 29 800 89 831
rect -89 -831 -29 -800
rect 29 -831 89 -800
rect -92 -847 -26 -831
rect -92 -881 -76 -847
rect -42 -881 -26 -847
rect -92 -897 -26 -881
rect 26 -847 92 -831
rect 26 -881 42 -847
rect 76 -881 92 -847
rect 26 -897 92 -881
<< polycont >>
rect -76 847 -42 881
rect 42 847 76 881
rect -76 -881 -42 -847
rect 42 -881 76 -847
<< locali >>
rect -263 1003 269 1013
rect -263 963 -255 1003
rect 255 963 269 1003
rect -263 959 -153 963
rect -249 949 -153 959
rect 153 959 269 963
rect 153 949 249 959
rect -249 887 -215 949
rect 215 887 249 949
rect -92 847 -76 881
rect -42 847 -26 881
rect 26 847 42 881
rect 76 847 92 881
rect -135 788 -101 804
rect -135 -804 -101 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 101 788 135 804
rect 101 -804 135 -788
rect -92 -881 -76 -847
rect -42 -881 -26 -847
rect 26 -881 42 -847
rect 76 -881 92 -847
rect -249 -949 -215 -887
rect 215 -949 249 -887
rect -249 -983 -153 -949
rect 153 -983 249 -949
rect -295 -2503 293 -2479
rect -295 -2543 -259 -2503
rect 251 -2543 293 -2503
rect -295 -2567 293 -2543
<< viali >>
rect -255 983 255 1003
rect -255 963 -153 983
rect -153 963 153 983
rect 153 963 255 983
rect -76 847 -42 881
rect 42 847 76 881
rect -135 -788 -101 788
rect -17 -788 17 788
rect 101 -788 135 788
rect -76 -881 -42 -847
rect 42 -881 76 -847
rect -259 -2543 251 -2503
<< metal1 >>
rect -99 881 -27 889
rect -99 847 -76 881
rect -42 847 -27 881
rect -99 843 -27 847
rect 25 881 97 889
rect 25 847 42 881
rect 76 847 97 881
rect 25 843 97 847
rect -88 841 -30 843
rect 30 841 88 843
rect -141 788 -95 800
rect -141 -788 -135 788
rect -101 -788 -95 788
rect -141 -800 -95 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 95 788 141 800
rect 95 -788 101 788
rect 135 -788 141 788
rect 95 -800 141 -788
rect -88 -847 -30 -841
rect -88 -881 -76 -847
rect -42 -881 -30 -847
rect -88 -887 -30 -881
rect 30 -847 88 -841
rect 30 -881 42 -847
rect 76 -881 88 -847
rect 30 -887 88 -881
rect -295 -2503 293 -2479
rect -295 -2543 -259 -2503
rect 251 -2543 293 -2503
rect -295 -2567 293 -2543
<< properties >>
string FIXED_BBOX -232 -966 232 966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 0.3 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
